-------------------------------------------------------------------------------
--
-- Title       : LL_SW_2_1_16_clk
-- Design      : 
-- Author      : Jean-Alexis Boulet
-- Company     : Telops
--
-------------------------------------------------------------------------------
--
-- Description : LocalLink Switch (mux) 2 to 1
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library Common_HDL;
use Common_HDL.Telops.all;

entity LL_SW_2_1_16_clk is 
   port(
      RX0_MOSI : in  t_ll_mosi;
      RX0_MISO : out t_ll_miso;
      
      RX1_MOSI : in  t_ll_mosi;
      RX1_MISO : out t_ll_miso;
      
      TX_MOSI  : out t_ll_mosi;
      TX_MISO  : in  t_ll_miso;
      
      SEL      : in  std_logic_vector(1 downto 0);
      
      ARESET      : in  std_logic;
      CLK         : in  STD_LOGIC
      );
end LL_SW_2_1_16_clk;


architecture RTL of LL_SW_2_1_16_clk is

signal RX_MOSI_DVAL_i : std_logic;
signal RX_MOSI_EOF_i : std_logic;
signal RX_MOSI_SOF_i : std_logic;
signal SEL_i     :std_logic_vector(1 downto 0);

begin    
   
   TX_MOSI.SUPPORT_BUSY <= '1';   
   
   SOF_sel : with SEL_i(0) select RX_MOSI_SOF_i <=
   RX0_MOSI.SOF when '0',   
   RX1_MOSI.SOF when others; 
   
   TX_MOSI.SOF <= RX_MOSI_SOF_i;

   EOF_sel : with SEL_i(0) select RX_MOSI_EOF_i <=
   RX0_MOSI.EOF when '0',   
   RX1_MOSI.EOF when others;
   
   TX_MOSI.EOF <= RX_MOSI_EOF_i;
     
   DATA_sel : with SEL_i(0) select TX_MOSI.DATA <= 
   RX0_MOSI.DATA when '0',
   RX1_MOSI.DATA when others;
      
   DVAL_sel : with SEL_i select RX_MOSI_DVAL_i <= 
   RX0_MOSI.DVAL when "00",   
   RX1_MOSI.DVAL when "01",
   '0'              when others;
   
   TX_MOSI.DVAL <= RX_MOSI_DVAL_i; 
  
   RX0_MISO.AFULL <= TX_MISO.AFULL;  
   RX1_MISO.AFULL <= TX_MISO.AFULL;   
   
   RX0_MISO.BUSY <= TX_MISO.BUSY when SEL_i = "00" else '1';         
   RX1_MISO.BUSY <= TX_MISO.BUSY when SEL_i = "01" else '1';
      
   ----------------------------------------------------------
   -- The classic switch
   ----------------------------------------------------------
   --SEL_i <= SEL; -- No change
  
   SEL_i <= "11" when ARESET = '1' else SEL; 
      
--   if ARESET = '1' then            
--      SEL_i <= "11"; -- Busy at reset                           
--   else
--      SEL_i <= SEL;
--   end if;
 
end RTL;
