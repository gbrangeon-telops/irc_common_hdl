------------------------------------------------------------------
--!   @file : mglk_DOUT_DVALiter
--!   @brief
--!   @details
--!
--!   $Rev$
--!   $Author$
--!   $Date$
--!   $Id$
--!   $URL$
------------------------------------------------------------------

-- ENO 27 sept 2017 :  
--    revision en profondeur pour tenir compte de le necessit� de sortir les donn�es hors AOI.
--    le flushing des fifos est abandonn�. le frame sync ne sert qu'� l'initialisation. Ainsi, le mode IWR sera facilit� puisque frame_sync est une entrave dans ce cas.  

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;
use work.fpa_define.all;
use work.fpa_common_pkg.all; 

entity afpa_lsync_mode_mux is
   port (
      ARESET          : in std_logic;
      CLK             : in std_logic;
      
      FPA_INTF_CFG    : in fpa_intf_cfg_type;
      
      READOUT_INFO_I  : in readout_info_type;
      READOUT_INFO_O  : out readout_info_type;
      
      LINE_GEN_ENABLE : out std_logic_vector(1 downto 0);
      
      READOUT         : in std_logic;
      DIN             : in std_logic_vector(57 downto 0);
      DIN_DVAL        : in std_logic
      
      );  
end afpa_lsync_mode_mux;


architecture rtl of afpa_lsync_mode_mux is
   
   component sync_reset
      port(
         ARESET : in std_logic;
         SRESET : out std_logic;
         CLK : in std_logic);
   end component;
   
   component double_sync is
      generic(
         INIT_VALUE : bit := '0'
         );
      port(
         D     : in std_logic;
         Q     : out std_logic := '0';
         RESET : in std_logic;
         CLK   : in std_logic
         );
   end component;
   
   type line_mux_fsm_type is (init_st1, init_st2, init_st3, init_st4, sync_flow_st);
   signal line_mux_fsm     : line_mux_fsm_type;
   signal sreset            : std_logic;
   signal pix_count         : unsigned(7 downto 0);   
   signal readout_info_pipe : readout_info_type;
   signal frame_sync        : std_logic;
   signal line_gen_enable_i : unsigned(1 downto 0);
   signal din_dval_i        : std_logic;
   signal sol_last          : std_logic;
   
   --attribute dont_touch     : string;
   --attribute dont_touch of dout_dval_o         : signal is "true"; 
   --attribute dont_touch of dout_o              : signal is "true";
   --attribute dont_touch of samp_fifo_ovfl      : signal is "true";
   --attribute dont_touch of flag_fifo_ovfl      : signal is "true";
   
begin
   
   --------------------------------------------------
   -- Outputs map
   -------------------------------------------------- 
   READOUT_INFO_O <= readout_info_pipe;
   LINE_GEN_ENABLE <= std_logic_vector(line_gen_enable_i);
   
   --------------------------------------------------
   -- synchro 
   --------------------------------------------------   
   U1A: sync_reset
   port map(
      ARESET => ARESET,
      CLK    => CLK,
      SRESET => sreset
      );      
   
   --------------------------------------------------
   -- Process
   --------------------------------------------------
   U2: process(CLK)
      variable incr :std_logic_vector(1 downto 0);
   begin
      if rising_edge(CLK) then         
         if sreset = '1' then      -- tant qu'on est en mode diag, la fsm est en reset.      
            line_mux_fsm <= init_st1;
            line_gen_enable_i <= (others => '0');
            -- pragma translate_off
            line_mux_fsm <= sync_flow_st;
            -- pragma translate_on
            
         else           
            
            frame_sync <= DIN(57);             -- sync_flag 
            din_dval_i <= DIN_DVAL;           
            
            readout_info_pipe <= READOUT_INFO_I;      -- delai requis pour une synchro avec line_gen_enable_i (tr�s important!)
            
            sol_last <= READOUT_INFO_I.SOL;
            
            case line_mux_fsm is         -- ENO: 23 juillet 2014. les etats init_st sont requis pour �viter des probl�mes de synchro          
               
               when init_st1 =>      
                  pix_count <= (others => '0');
                  if frame_sync = '1' then  -- je vois un signal de synchro
                     line_mux_fsm <= init_st2;
                  end if;                                                                       
               
               when init_st2 =>     
                  if frame_sync = '0' then  -- je ne vois plus le signal de synchro
                     line_mux_fsm <= init_st3;
                  end if;  
               
               when init_st3 =>
                  if din_dval_i = '1' then      
                     pix_count <= pix_count + DEFINE_FPA_TAP_NUMBER;
                  end if;                                           
                  if pix_count >= 64 then    -- je vois au moins un nombre de pixels �quivalent � la plus petite ligne d'image de TEL-2000. cela implique que le syst�me en amont est actif. je m'en vais en idle et attend la prochaine synchro 
                     line_mux_fsm <= init_st4;     
                  end if;
               
               when init_st4 =>             -- la carte ADc est connect�e sinon on ne parviendra pas ici
                  if READOUT_INFO_I.READ_END = '1' then  -- je vois la tomb�e du fval d'une readout_info =>
                     line_mux_fsm <= sync_flow_st; 
                  end if;
                  
               -- une fois ici, je suis certain que les deux flows seront synchronisables
               when sync_flow_st =>
                  if READOUT_INFO_I.SOL = '1' and sol_last = '0' then 
                     line_gen_enable_i <= not line_gen_enable_i; -- on commute indefininement entre les synchronisateurs de lignes
                  end if;
                                 
               when others =>
               
            end case;
            
         end if;
      end if;
   end process;
   
end rtl;