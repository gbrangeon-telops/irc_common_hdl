------------------------------------------------------------------
--!   @file fpa_intf_sequencer
--!   @brief sequenceur du modeule FPA interface
--!   @details ce module assure la coordination des activit�s dans le module FPA Interface
--! 
--!   $Rev$
--!   $Author$
--!   $Date$
--!   $Id$
--!   $URL$
------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all; 
use work.fpa_common_pkg.all;        -- pour connaitre le type d'interface du projet
use work.FPA_Define.all;
use work.Proxy_Define.all;

entity fpa_intf_sequencer is
   
   generic (       
      BYPASS_FPA_PROTECTION : boolean := false  -- en simulation, permet de contourner  toutes les protections. Doit toujours d�meurer � false en mode r�el 
      );
   
   port(       
      --------------------------------------------------
      -- INPUTS
      --------------------------------------------------
      CLK                : in std_logic;
      ARESET             : in std_logic;       
      FPA_INTF_CFG       : in fpa_intf_cfg_type; --! configuration           
      TRIG_CTLER_STAT    : in std_logic_vector(7 downto 0); --! statuts du gestionnaire des trigs du FPA          
      FPA_DRIVER_STAT    : in std_logic_vector(31 downto 0); --! statuts du pilote Hardware du FPA     
      FPA_COOLER_STAT    : in fpa_cooler_stat_type; --! statut du refroidisseur     
      FPA_HARDW_STAT     : in fpa_hardw_stat_type; --! statut (type + mise-�-jour) de toutes les cartes de proximit� (proxy, flex, DDC, ADC, harnais etc...)   
      FPA_SOFTW_STAT     : in fpa_firmw_stat_type;--
      FPA_VHD_STAT       : in fpa_firmw_stat_type;--
      FPA_TEMP_STAT      : in fpa_temp_stat_type; --! statut du lecteur de temp�rature
      --------------------------------------------------
      -- OUTPUTS
      --------------------------------------------------     
      TRIG_CTLER_EN      : out std_logic; --! controle du gestionnaire des trigs      
      FPA_DRIVER_EN      : out std_logic; --! controle du pilote Hardware du FPA      
      FPA_POWER          : out std_logic; --! controle de l'allumage du FPA    
      INTF_SEQ_STAT      : out std_logic_vector(7 downto 0); --! statut du s�quenceur     
      DIAG_MODE_ONLY     : out std_logic  --! diag mode only. � '1' <=> seul le mode diag est autoris�      
      );
end fpa_intf_sequencer;



architecture RTL of fpa_intf_sequencer is  
   
   component sync_reset
      port(
         ARESET : in STD_LOGIC;
         SRESET : out STD_LOGIC;
         CLK    : in STD_LOGIC);
   end component;
   
   component Clk_Divider is
      Generic(	Factor:		integer := 2);		
      Port ( Clock  : in std_logic;
         Reset  : in std_logic;		
         Clk_div: out std_logic);
   end component;
   
   type status_type is (not_available, success, failure);
   type fpa_sequencer_sm_type is (init_st1, init_st2, idle, trig_ctrl_st, active_prog_st, wait_trig_done_st, wait_prog_end_st, trig_en_st);
   signal fpa_hardw_up2date   : status_type;
   signal fpa_hardw_type      : status_type;
   signal fpa_vhd_stat_i      : status_type;
   signal fpa_softw_stat_i    : status_type;
   signal fpa_temp_stat_i     : status_type;
   signal hardw_global_status : status_type;
   signal firmw_global_status : status_type;
   signal fpa_sequencer_sm    : fpa_sequencer_sm_type;
   signal sreset              : std_logic;
   --signal fpa_intf_type_err_i : std_logic;
   signal fpa_power_i           : std_logic;
   signal trig_ctler_en_i     : std_logic; 
   signal fpa_driver_en_i     : std_logic;
   signal trig_ctler_done     : std_logic;
   signal fpa_driver_done     : std_logic;
   signal fpa_driver_rqst     : std_logic; -- permet de saboir si le pilote hw requiert de reprogrammer le FPA
   signal fpa_cooler_on       : std_logic;
   signal done                : std_logic; 
   signal fpa_hardw_err       : std_logic;
   signal diag_mode_only_i    : std_logic;
   signal fpa_softw_err       : std_logic;
   signal fpa_vhd_err         : std_logic;
   signal fpa_init_cfg_rdy    : std_logic;
   
   
   
   --   attribute keep : string;
   --   attribute keep of CLK_1sec : signal is "true";
   
begin    
   
   
   --------------------------------------------------
   -- mapping des sorties
   -------------------------------------------------- 
   FPA_POWER <= fpa_power_i;
   TRIG_CTLER_EN <= trig_ctler_en_i;
   FPA_DRIVER_EN <= fpa_driver_en_i;
   DIAG_MODE_ONLY <= diag_mode_only_i;
   
   --stat                     
   INTF_SEQ_STAT(7 downto 4) <= (others => '0');   
   INTF_SEQ_STAT(3) <= fpa_softw_err; 
   INTF_SEQ_STAT(2) <= fpa_vhd_err; 
   INTF_SEQ_STAT(1) <= fpa_hardw_err;           
   INTF_SEQ_STAT(0) <= done; 
   
   --------------------------------------------------
   -- mapping des entrees
   -------------------------------------------------- 
   fpa_driver_rqst <= FPA_DRIVER_STAT(1);
   trig_ctler_done <= TRIG_CTLER_STAT(0);
   fpa_driver_done <= FPA_DRIVER_STAT(0);   
   
   --------------------------------------------------
   -- Sync reset
   -------------------------------------------------- 
   U1 : sync_reset
   port map(ARESET => ARESET, CLK => CLK, SRESET => sreset); 
   
   -----------------------------------------------------------
   -- V�rification des statuts des cartes �lectroniques 
   -----------------------------------------------------------
   U2: process(CLK)
   begin          
      if rising_edge(CLK) then         
         
         if FPA_HARDW_STAT.DVAL = '1' and FPA_VHD_STAT.DVAL = '1' then     -- dval est requis pour eviter de sortir des fausses erreurs
            
            -- on v�rifie que le montage �lectronique est conforme au design vhd et on v�rifie aussi que les IO de contr�le du FPGA sont conformes aux specs de l'iDDCA
            if FPA_HARDW_STAT.IDDCA_INFO.FPA_ROIC = FPA_VHD_STAT.FPA_ROIC and  FPA_HARDW_STAT.IDDCA_INFO.FPA_OUTPUT = FPA_VHD_STAT.FPA_OUTPUT and  FPA_HARDW_STAT.IDDCA_INFO.FPA_INPUT = FPA_VHD_STAT.FPA_INPUT then  -- FPA_VHD_STAT.FPA_ROIC est une reference s�re car cod� en hardware.              
               fpa_hardw_type <= success;                                                                                                                                                                       ---- FPA_HARDW_STAT.IDDCA_INFO.FPA_INPUT provient des cartes d'interface des d�tecteurs et FPA_VHD_STAT.FPA_INPUT provient d'un module qui mesure la tension du FPGA          
               fpa_hardw_err <= '0';
            else
               fpa_hardw_type <= failure;
               fpa_hardw_err <= '1';
            end if; 
            
            -- on v�rifie que l'�lectronique est � jour
            -- if FPA_HARDW_STAT.HARDW_UP2DATE = '1' then
            fpa_hardw_up2date <= success;
            --   fpa_hardw_err <= '0';
            --else
            --   fpa_hardw_up2date <= failure;
            --   fpa_hardw_err <= '1';
            --end if;
            
         else                
            fpa_hardw_up2date <= not_available;
            fpa_hardw_type <= not_available;
            fpa_hardw_err <= '0';            
         end if;
         
      end if;
   end process; 
   
   -----------------------------------------------------------
   -- V�rification des statuts du firmware 
   -----------------------------------------------------------
   U3: process(CLK)
   begin          
      if rising_edge(CLK) then 
         if sreset = '1' then 
            fpa_vhd_stat_i <= not_available; 
            fpa_softw_stat_i <= not_available;
            fpa_vhd_err <= '0';
            fpa_softw_err <= '0';
         else
            
            -- on v�rifie que le design Vhd est conforme � FPA_define(Ceci est requis car tous les defines ont le m�me nom)
            if FPA_VHD_STAT.DVAL = '1' then               
               if FPA_VHD_STAT.FPA_ROIC = DEFINE_FPA_ROIC and FPA_VHD_STAT.FPA_OUTPUT = DEFINE_FPA_OUTPUT then  
                  fpa_vhd_stat_i <= success;
                  fpa_vhd_err <= '0';
               else
                  fpa_vhd_stat_i <= failure;
                  fpa_vhd_err <= '1';
               end if;
            else
               fpa_vhd_stat_i <= not_available;
               fpa_vhd_err <= '0';
            end if;
            --
            -- on v�rifie que les pilotes software (PPC/�Blaze) sont conformes � la definition dans FPA_define
            if FPA_SOFTW_STAT.DVAL = '1' then           -- dval est requis car cela prend du temps au PPC pour envoyer l'info au Hardw
               if FPA_SOFTW_STAT.FPA_ROIC = DEFINE_FPA_ROIC and FPA_SOFTW_STAT.FPA_OUTPUT = DEFINE_FPA_OUTPUT then 
                  fpa_softw_stat_i <= success;
                  fpa_softw_err <= '0';
               else
                  fpa_softw_stat_i <= failure;
                  fpa_softw_err <= '1';
               end if;
            else
               fpa_softw_stat_i <= not_available;  --! requis car il y a un delai avant que l'init de PPC envoie cette information
               fpa_softw_err <= '0';
            end if;
            -- 
         end if;
      end if;
   end process; 
   
   -----------------------------------------------------------
   -- V�rification du statut du refroidisseur de la cfg d'initisalisation
   -----------------------------------------------------------
   -- on v�rifie que le refroidisseur est allum� 
   -- on v�rifie que la config d'initialisation est pr�te
   U5: process(CLK)
   begin          
      if rising_edge(CLK) then 
         fpa_cooler_on <= FPA_COOLER_STAT.COOLER_ON;
         fpa_init_cfg_rdy <= (DEFINE_FPA_INIT_CFG_NEEDED and FPA_INTF_CFG.COMN.FPA_INIT_CFG_RECEIVED) or not DEFINE_FPA_INIT_CFG_NEEDED; 
      end if;
   end process;  
   
   -----------------------------------------------------------
   -- V�rification de la temperature du d�tecteur  
   -----------------------------------------------------------
   -- on v�rifie que la temp�rature lue est conforme pour 
   -- l'allumage du d�tecteur
   U6: process(CLK)
   begin          
      if rising_edge(CLK) then 
         if FPA_TEMP_STAT.FPA_PWR_ON_TEMP_REACHED = '1' then
            fpa_temp_stat_i <= success;
         else
            fpa_temp_stat_i <= failure;
         end if;
         
         -- pragma translate_off
         if BYPASS_FPA_PROTECTION = true then
            fpa_temp_stat_i <= success;
         end if;         
         -- pragma translate_on
         
      end if;
   end process;
   
   -----------------------------------------------------------
   -- Compilation des diff�rents statuts pr�-allumage  
   -----------------------------------------------------------
   -- on compile les diff�rents statuts p�-allumage 
   U7: process(CLK)
   begin          
      if rising_edge(CLK) then
         
         -- compilation des statuts du hw (type de cartes et mises-�-jour)
         if fpa_hardw_up2date = not_available or fpa_hardw_type = not_available then
            hardw_global_status <= not_available;
         elsif fpa_hardw_up2date = success and fpa_hardw_type = success then
            hardw_global_status <= success;
         else
            hardw_global_status <= failure;
         end if;
         
         -- pragma translate_off
         if BYPASS_FPA_PROTECTION = true then
            hardw_global_status <= success;
         end if;         
         -- pragma translate_on
         
         -- compilation des statuts firmware (vhd et du software (PPC/�Blaze))
         if fpa_softw_stat_i = not_available or fpa_vhd_stat_i = not_available then 
            firmw_global_status <= not_available;
         elsif fpa_softw_stat_i = success and fpa_vhd_stat_i = success then 
            firmw_global_status <= success;                                
         else
            firmw_global_status <= failure;
         end if;
         
         -- pragma translate_off
         if BYPASS_FPA_PROTECTION = true then
            firmw_global_status <= success;
         end if;         
         -- pragma translate_on
         
      end if;      
   end process;     
   
   --------------------------------------------------
   -- Allumage du Flex ou du Proxy  
   -------------------------------------------------- 
   -- il faut que ce soit un process totalement ind�pendant qui 
   -- s'occupe de l'allumage des cartes sensibles
   U8: process(CLK)
   begin          
      if rising_edge(CLK) then 
         if sreset = '1' then 
            fpa_power_i <= '0'; 
         else                      
            -- le proxy ou le FPA ne peut s'allumer que ssi : 
            -- 1) le hawdware et le firmare sont conformes
            -- 2) le refroidisseur est en fonction
            -- 3) la temp�rature du d�tecteur est conforme
            -- 4) on re�oit l'ordre d'allumage en provenance du PPC/�Blaze
            -- 5) le statut relatif � la config d'initialisation est conforme
            if hardw_global_status = success and firmw_global_status = success and fpa_temp_stat_i = success then 
               fpa_power_i <= FPA_INTF_CFG.COMN.FPA_PWR_ON and fpa_cooler_on and fpa_init_cfg_rdy; 
            else
               fpa_power_i <= '0';
            end if;            
         end if;
      end if;
   end process;    
   
   --------------------------------------------------
   -- sequenceur
   --------------------------------------------------   
   --
   U9: process(CLK)
   begin          
      if rising_edge(CLK) then 
         if sreset = '1' then 
            fpa_sequencer_sm <= init_st1;
            trig_ctler_en_i <= '0';
            fpa_driver_en_i <= '0';
            done <= '0';
            diag_mode_only_i <= '0'; 
            
         else             
            
            case fpa_sequencer_sm is 
               
               when init_st1 => 
                  done <= '0';
                  trig_ctler_en_i <= '0';
                  fpa_driver_en_i <= '0';
                  diag_mode_only_i <= '0'; 
                  if firmw_global_status = success then 
                     fpa_sequencer_sm <= init_st2; 
                  else     -- statut non encore disponible ou failure, rien � faire sauf attendre
                  end if;
               
               when init_st2 =>
                  diag_mode_only_i <= '1'; -- si le firmware est correct, au moins le mode diag est possible. 
                  if hardw_global_status = success then                        
                     fpa_sequencer_sm <= idle;
                  elsif hardw_global_status = failure then     
                     fpa_sequencer_sm <= idle;
                  else  -- statut non encore disponible, on attend
                     trig_ctler_en_i <= FPA_INTF_CFG.COMN.FPA_DIAG_MODE; -- le contr�leur de trig est activ� si le mode diag est demand�. Sinon , rien ne se passe
                  end if;                  
               
               when idle =>      -- on ne vient ici que lorsqu'au moins le firmware est correct                    
                  done <= '1';
                  if diag_mode_only_i = '1' then   
                     trig_ctler_en_i <= FPA_INTF_CFG.COMN.FPA_DIAG_MODE; -- en mode diag_only le contr�leur de trigs est en fonction ssi le mode diag est demand�.
                  end if;                  
                  if fpa_power_i = '1' then      -- certes fpa_power_i est l'ordre d'allumage mais ne dit pas si le fpa est allum� r�ellement ou pas. Mais ce n'est pas grave car fpa �teint => fpa_driver_rqst = '0'
                     diag_mode_only_i <= '0';    -- le mode diag n'est plus le seul mode une fois que le d�tecteur est allum�
                     if fpa_driver_rqst = '1' then 
                        fpa_sequencer_sm <= trig_ctrl_st;
                     end if;
                  else                         
                     diag_mode_only_i <= '1';   -- le mode diag uniquement si le d�tecteur n'est pas encore allum� (cooldown ou pas d'ordre d'allumage)
                  end if;                    
               
               when trig_ctrl_st =>  -- si on vient ici, c'est que le d�tecteur est allum� et qu'on veuille le programmer
                  if PROG_FREE_RUNNING_TRIG = '1' then   -- en mode free_running_trig, il n'est pas necessaire d'arr�ter le contr�leur de trig avant programmation
                     fpa_sequencer_sm <= active_prog_st;
                     trig_ctler_en_i <= '1';  -- on s'assure que les trigs sont envoy�s au d�tecteur avant de le programmer (cas des scd par exemple)
                  else                     
                     fpa_sequencer_sm <= wait_trig_done_st;
                     trig_ctler_en_i <= '0'; -- on arrete tout trig avant de programmer le d�tecteur (cas de plusieurs d�tecteurs analogiques)
                  end if;
               
               when wait_trig_done_st =>    
                  if trig_ctler_done = '1' then 
                     fpa_sequencer_sm <= active_prog_st;
                  end if;
               
               when active_prog_st =>                -- on programme le FPA
                  fpa_driver_en_i <= '1';
                  if fpa_driver_done = '0' then 
                     fpa_sequencer_sm <= wait_prog_end_st;
                  end if;    
               
               when wait_prog_end_st =>        -- on attend la fin de la programmation                
                  fpa_driver_en_i <= '0';    
                  if fpa_driver_done = '1' then 
                     fpa_sequencer_sm <= trig_en_st;
                  end if; 
               
               when trig_en_st =>            -- on permet les integrations 
                  trig_ctler_en_i <= '1';
                  fpa_sequencer_sm <= idle; 
               
               when others =>
               
            end case;      
            
         end if;
      end if;
   end process;
   
end RTL;
