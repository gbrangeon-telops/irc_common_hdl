---------------------------------------------------------------------------------------------------
--                                                      ..`??!````??!..
--                                                  .?!                `1.
--                                               .?`                      i
--                                             .!      ..vY=!``?74.        i
--.........          .......          ...     ?      .Y=` .+wA..   ?,      .....              ...
--"""HMM"""^         MM#"""5         .MM|    :     .H\ .JQgNa,.4o.  j      MM#"MMN,        .MM#"WMF
--   JM#             MMNggg2         .MM|   `      P.;,jMt   `N.r1. ``     MMmJgMM'        .MMMNa,.
--   JM#             MM%````         .MM|   :     .| 1A Wm...JMy!.|.t     .MMF!!`           . `7HMN
--   JMM             MMMMMMM         .MMMMMMM!     W. `U,.?4kZ=  .y^     .!MMt              YMMMMB=
--                                          `.      7&.  ?1+...JY'     J
--                                           ?.        ?""""7`       .?`
--                                             :.                ..?`
--                                               `!...........??`
---------------------------------------------------------------------------------------------------
--
-- Title       : LocalLink_Fifo
-- Design      : VP30
-- Author      : Patrick Daraiche
-- Company     : Telops Inc.
--
--  $Revision: 
--  $Author: 
--  $LastChangedDate:
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;    
use work.fpa_common_pkg.all;

entity LL8_ext_fifo8 is
   generic(
      FifoSize		   : integer := 256;  -- 256
      Latency        : integer := 32;  -- Input module latency (to control RX_LL_MISO.AFULL)      
      ASYNC          : boolean := true);	-- Use asynchronous fifos
   port(
      --------------------------------
      -- FIFO RX Interface
      --------------------------------
      RX_LL_MOSI  : in  t_ll_ext_mosi8;
      RX_LL_MISO  : out t_ll_ext_miso;
      CLK_RX 		: in 	std_logic;
      FULL        : out std_logic;
      WR_ERR      : out std_logic;
      --------------------------------
      -- FIFO TX Interface
      --------------------------------
      TX_LL_MOSI  : out t_ll_ext_mosi8;
      TX_LL_MISO  : in  t_ll_ext_miso;
      CLK_TX 		: in 	std_logic;
      EMPTY       : out std_logic; -- This signal should actually be called "IDLE"
      --------------------------------
      -- Common Interface
      --------------------------------
      ARESET		: in std_logic
      );
end LL8_ext_fifo8;

architecture RTL of LL8_ext_fifo8 is 
   
   component sync_reset
      port(
         ARESET : in std_logic;
         SRESET : out std_logic;
         CLK : in std_logic);
   end component;
   
   component sfifo_w10_d256
      port(
         clk : in std_logic;
         din : in std_logic_vector(9 downto 0);
         rd_en : in std_logic;
         srst : in std_logic;
         wr_en : in std_logic;
         data_count : out std_logic_vector(7 downto 0);
         dout : out std_logic_vector(9 downto 0);
         empty : out std_logic;
         full : out std_logic;
         overflow : out std_logic;
         valid : out std_logic);
   end component;  
   
   signal fifo_count_256  : std_logic_vector(7 downto 0);   
   signal fifo_dout : std_logic_vector(9 downto 0);
   signal fifo_din : std_logic_vector(9 downto 0);
   signal fifo_rd_ack : std_logic;			
   signal fifo_rd_en : std_logic;
   
   signal hold_dval  : std_logic;
   signal TX_DVAL_buf: std_logic;
   signal FULLi      : std_logic;    
   signal AFULLi     : std_logic;    
   signal WR_ERRi    : std_logic;
   signal EMPTYi     : std_logic;
   signal fifo_wr_en : std_logic;
   
   signal FoundGenCase : boolean;      
   signal RESET_TX : std_logic;                  
   signal RESET_RX : std_logic;   
   
   -- This signal is for debug only and will be optimized out by xst
   signal tx_cnt     : unsigned(31 downto 0); 
   --   attribute keep    : string; 
   --   attribute keep of tx_cnt : signal is "true";     
   
begin      
   
   sync_RESET_TX :  sync_reset
   port map(ARESET => ARESET, SRESET => RESET_TX, CLK => CLK_TX); 
   
   sync_RESET_RX :  sync_reset
   port map(ARESET => ARESET, SRESET => RESET_RX, CLK => CLK_RX);
   
      
   gen_8_256 : if (FifoSize > 32 and FifoSize <= 256 and not ASYNC) generate
      begin
      FoundGenCase <= true;
      AFULLi <= '1' when (unsigned(fifo_count_256) > (255-(Latency+1)) or FULLi = '1') else '0';
      sfifo_w10_d256_inst : sfifo_w10_d256
      port map(
         clk => CLK_RX,
         din => fifo_din,
         rd_en => fifo_rd_en,
         srst => RESET_TX,
         wr_en => fifo_wr_en,
         data_count => fifo_count_256,
         dout => fifo_dout,
         empty => EMPTYi,
         full => FULLi,
         overflow => WR_ERRi,
         valid => fifo_rd_ack
         );
   end generate gen_8_256;	
   
   
   TX_LL_MOSI.SUPPORT_BUSY <= '1';
   
   -- Fifo write control
   fifo_wr_en <= RX_LL_MOSI.DVAL and not FULLi;
   
   -- Fifo read control
   fifo_rd_en <= not TX_LL_MISO.AFULL and not (TX_LL_MISO.BUSY and TX_DVAL_buf);
   
   -- Write interface signals
   fifo_din <= (RX_LL_MOSI.SOF & RX_LL_MOSI.EOF & RX_LL_MOSI.DATA);	
   
   -- OUTPUT MAPPING                       
   TX_LL_MOSI.DVAL <= TX_DVAL_buf when FoundGenCase else '0';
   TX_DVAL_buf <= fifo_rd_ack or hold_dval;
   TX_LL_MOSI.DATA <= fifo_dout(7 downto 0) when FoundGenCase else (others => '0');
   TX_LL_MOSI.EOF <= fifo_dout(8) when FoundGenCase else '0';	 
   TX_LL_MOSI.SOF <= fifo_dout(9) when FoundGenCase else '0';                  
   
   FULL <= FULLi when FoundGenCase else '1'; 
   --RX_LL_MISO.AFULL <= AFULLi when FoundGenCase else '1'; 
   
   no_latency : if Latency = 0 generate
      RX_LL_MISO.AFULL <= '0';
   end generate no_latency;        
   
   with_latency : if Latency > 0 generate   
      -- PDU: We register AFULL to help timing closure. Anyway one extra clock cycle on 
      -- AFULL should not matter in the vast majority of cases. Just to make sure, we
      -- added +1 to the generic Latency.
      process (CLK_RX)
      begin                  
         if rising_edge(CLK_RX) then      
            if FoundGenCase then
               RX_LL_MISO.AFULL <= AFULLi or RESET_RX;
            else
               RX_LL_MISO.AFULL <= '1';   
            end if;    
         end if;
      end process;
   end generate with_latency;      
   
   
   RX_LL_MISO.BUSY <= FULLi or RESET_RX;
   WR_ERR <= WR_ERRi when FoundGenCase else '0'; 
   
   -- DVALID latch (when RX is not ready, all we have to do is hold the DVal signal, the fifo interface does the rest)
   tx_proc : process (CLK_TX)
   begin	
      if rising_edge(CLK_TX) then
         if RESET_TX = '1' then
            hold_dval <= '0';
            tx_cnt <= (others => '0');
         else
            if TX_DVAL_buf = '1' and TX_LL_MISO.BUSY = '0' then
               tx_cnt <= tx_cnt + 1;
            end if;
            
            hold_dval <= TX_LL_MISO.BUSY and TX_DVAL_buf;  
            -- pragma translate_off   
            assert (FoundGenCase or FifoSize = 0) report "Invalid LocalLink fifo generic settings!" severity FAILURE;
            if FoundGenCase then
               assert (WR_ERRi /= '1') report "LocalLink fifo overflow!!!" severity ERROR;
            end if;
            -- pragma translate_on
         end if;		
      end if;
   end process;   
   
   rx_proc : process (CLK_RX)
      variable empty_mid : std_logic;
   begin	
      if rising_edge(CLK_RX) then
         if RESET_RX = '1' or EMPTYi = '0' or TX_DVAL_buf = '1' then
            empty_mid := '0';
            EMPTY <= '0';
         else
            empty_mid := EMPTYi;
            EMPTY <= empty_mid;
         end if;		
      end if;
   end process;
   
end RTL;
