-------------------------------------------------------------------------------
--
--      Project:  Aurora Module Generator
--
--         Date:  $Date$
--          Tag:  $Name: i+IP+125372 $
--         File:  $RCSfile: sim_reset_on_configuration_vhd.ejava,v $
--          Rev:  $Revision$
--
--      Company:  Xilinx
-- Contributors:  R. K. Awalt, B. L. Woodard, N. Gulstone, N. Jayarajan
--
--   Disclaimer:  XILINX IS PROVIDING THIS DESIGN, CODE, OR
--                INFORMATION "AS IS" SOLELY FOR USE IN DEVELOPING
--                PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY
--                PROVIDING THIS DESIGN, CODE, OR INFORMATION AS
--                ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE,
--                APPLICATION OR STANDARD, XILINX IS MAKING NO
--                REPRESENTATION THAT THIS IMPLEMENTATION IS FREE
--                FROM ANY CLAIMS OF INFRINGEMENT, AND YOU ARE
--                RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY
--                REQUIRE FOR YOUR IMPLEMENTATION.  XILINX
--                EXPRESSLY DISCLAIMS ANY WARRANTY WHATSOEVER WITH
--                RESPECT TO THE ADEQUACY OF THE IMPLEMENTATION,
--                INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR
--                REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE
--                FROM CLAIMS OF INFRINGEMENT, IMPLIED WARRANTIES
--                OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
--                PURPOSE.
--
--                (c) Copyright 2004 Xilinx, Inc.
--                All rights reserved.
--

--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--   __  __ 
--  /   /\/   / 
-- /__/  \  /    Vendor: Xilinx 
-- \   \   \/     Version : 1.0
--  \   \         Application : RocketIO Wizard 
--  /   /         Filename : mgt_wrapper.vhd
-- /__/   /\     Timestamp : 02/08/2005 09:12:43
-- \   \  /  \ 
--  \__\/\__\ 
--
--
-- Module MGT_WRAPPER 
-- Generated by Xilinx RocketIO Wizard, generation mechanism modified for COREGen Aurora

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- synopsys translate_off
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
-- synopsys translate_on

--***************************** Entity Declaration *****************************
entity aurora_sim_reset_on_config is
port 
(
    GSR_IN     : in std_logic
);
end aurora_sim_reset_on_config;

architecture BEHAVIORAL of aurora_sim_reset_on_config is
  
-- translate_off
    component ROCBUF 
    port 
    ( 
        I : in std_logic; 
        O : out std_logic 
    ); 
    end component; 
-- translate_on    

signal dummy_signal : std_logic;

                       

--********************************* Main Body of Code****************************
                       
begin                      
-- translate_off   
    GSR <= GSR_IN;                       
    ------------------------------  ROCBUF Instantiation -----------------------   
    -- This component is required for correctly resetting the GT11 component on configuration
    -- It is for simulation alone and will be ripped out during synthesis.
    U1 : ROCBUF 
    port map 
    (
        I => GSR,
        O => open
    );               
-- translate_on  

  -- This code is useless but prevents XST from creating a blackbox.
  dummy_signal <= GSR_IN;


end BEHAVIORAL;
