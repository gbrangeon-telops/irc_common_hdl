---------------------------------------------------------------------------------------------------
--                                                      ..`??!````??!..
--                                                  .?!                `1.
--                                               .?`                      i
--                                             .!      ..vY=!``?74.        i
--.........          .......          ...     ?      .Y=` .+wA..   ?,      .....              ...
--"""HMM"""^         MM#"""5         .MM|    :     .H\ .JQgNa,.4o.  j      MM#"MMN,        .MM#"WMF
--   JM#             MMNggg2         .MM|   `      P.;,jMt   `N.r1. ``     MMmJgMM'        .MMMNa,.
--   JM#             MM%````         .MM|   :     .| 1A Wm...JMy!.|.t     .MMF!!`           . `7HMN
--   JMM             MMMMMMM         .MMMMMMM!     W. `U,.?4kZ=  .y^     .!MMt              YMMMMB=
--                                          `.      7&.  ?1+...JY'     .J
--                                           ?.        ?""""7`       .?`
--                                             :.                ..?`
--
---------------------------------------------------------------------------------------------------
--
-- Title       : DPB_Define
-- Design      : DPB (Data Processing Board)
-- Author      : Patrick Dubois
-- Company     : Telops Inc.
--
---------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library Common_HDL;
use Common_HDL.Telops.all;
use work.CAMEL_Define.all;

package DPB_Define is
   ------------------------------------------
   -- Constants
   ------------------------------------------
   constant CLINK_VERSION  : std_logic_vector(7 downto 0) := "110" & "00000";
   constant CLINK_HDR_VERSION: std_logic_vector(3 downto 0) := x"4";    -- default to version 3 header
   constant AMAX : integer := 26; -- DDR address space: 26 downto 0
   constant CACHE_INIT_PHASE : integer := -102;    
   
   constant INACTIVE_WB : t_wb_mosi := (x"0000", '0', x"000", '0', '0'); 
   
   -- Define number of bits used
   constant MAXFFTLEN: integer := 16;
   constant IMGLEN   : integer := 20;
   constant XLEN     : integer := 10;
   constant YLEN     : integer := 10;
   constant ZLEN     : integer := 24;
   constant PLLEN    : integer := 24;
   constant TAGLEN   : integer := 8;
   constant AVGLEN   : integer := 6;
   constant DIAGLEN  : integer := 16;
   constant LVALLEN  : integer := 16;
   constant FVALLEN  : integer := 16;
   constant HEADERLEN: integer := 16;
   constant LPAUSELEN: integer := 16;
   constant SBANDLEN : integer := MAXFFTLEN;
   constant PAGELEN  : integer := 22;
   constant DUILEN   : integer := 29;   
   constant DPBSTATLEN : integer := 64;
   constant PPCSTATLEN : integer := 16;
   constant CLINKMODELEN     : integer := 6;
   constant FRAMESPERCUBELEN : integer := 16;
   constant DIAGSIZELEN      : integer := 16;
   constant ACQNUMLEN        : integer := 10;
   constant DIAGMODELEN      : integer := 4;
   constant DPMODELEN        : integer := 8;
   constant DIAGROMLEN       : integer := 1024;
   
   constant BSQ : std_logic_vector(1 downto 0) := "00";
   constant BIP : std_logic_vector(1 downto 0) := "01";
   
   -- Data Processing Modes (8-bit). If MSB is '1', data is generated by pattern generator (diag mode).
   constant DP_STOP           : std_logic_vector(DPMODELEN-1 downto 0) := x"00";
   constant DP_IGM            : std_logic_vector(DPMODELEN-1 downto 0) := x"01";
   constant DP_RAW_SPC        : std_logic_vector(DPMODELEN-1 downto 0) := x"02";
   constant DP_CAL_SPC_ONLY   : std_logic_vector(DPMODELEN-1 downto 0) := x"03";
   constant DP_CAL_SPC_N_IGM  : std_logic_vector(DPMODELEN-1 downto 0) := x"04";
   constant DP_GAIN_OFFSET    : std_logic_vector(DPMODELEN-1 downto 0) := x"05";
   constant DP_HOT_BB_STORE   : std_logic_vector(DPMODELEN-1 downto 0) := x"06";
   constant DP_HOT_BB_OUT     : std_logic_vector(DPMODELEN-1 downto 0) := x"07";
   constant DP_COLD_BB_STORE  : std_logic_vector(DPMODELEN-1 downto 0) := x"08";
   constant DP_COLD_BB_OUT    : std_logic_vector(DPMODELEN-1 downto 0) := x"09";
   constant DP_RAW_SPC_N_IGM  : std_logic_vector(DPMODELEN-1 downto 0) := x"0A";
   constant DP_CAMERA         : std_logic_vector(DPMODELEN-1 downto 0) := x"0F";
   
   constant DP_DIAG_STOP           : std_logic_vector(DPMODELEN-1 downto 0) := x"80";
   constant DP_DIAG_IGM            : std_logic_vector(DPMODELEN-1 downto 0) := x"81";
   constant DP_DIAG_RAW_SPC        : std_logic_vector(DPMODELEN-1 downto 0) := x"82";
   constant DP_DIAG_CAL_SPC_ONLY   : std_logic_vector(DPMODELEN-1 downto 0) := x"83";
   constant DP_DIAG_CAL_SPC_N_IGM  : std_logic_vector(DPMODELEN-1 downto 0) := x"84";
   constant DP_DIAG_GAIN_OFFSET    : std_logic_vector(DPMODELEN-1 downto 0) := x"85";
   constant DP_DIAG_HOT_BB_STORE   : std_logic_vector(DPMODELEN-1 downto 0) := x"86";
   constant DP_DIAG_HOT_BB_OUT     : std_logic_vector(DPMODELEN-1 downto 0) := x"87";
   constant DP_DIAG_COLD_BB_STORE  : std_logic_vector(DPMODELEN-1 downto 0) := x"88";
   constant DP_DIAG_COLD_BB_OUT    : std_logic_vector(DPMODELEN-1 downto 0) := x"89";
   constant DP_DIAG_RAW_SPC_N_IGM  : std_logic_vector(DPMODELEN-1 downto 0) := x"8A";
   constant DP_DIAG_CAMERA         : std_logic_vector(DPMODELEN-1 downto 0) := x"8F";
   
   -- CameraLink Mode Settings (Are now bit positions for enabling features)
   constant CL_FULL_BIT  : integer := 0; -- Cameralink BASE_bar/FULL Mode selection bit position
   constant CL_LOOP_BIT  : integer := 1; -- Cameralink Internal LOOPBACK test bit position
   constant CL_RIOTX_BIT : integer := 2; -- Cameralink Transmit on RIO for external loopback bit position
   constant CL_DUAL_BIT  : integer := 3; -- Cameralink Enable DUAL ports in Base mode bit position
   constant CL_SWAP_BIT  : integer := 4; -- Cameralink Enable Pixel Byte Swapping (Pixel Endianness for Bitflow Board)
   constant CL_DATASWAP_BIT  : integer := 5; -- Cameralink Enable Pixel Byte Swapping for data only (Pixel Endianness for data part only)
   
   -- Reintroduced these constants, it doesn't hurt anyone ;)
   constant CLINK_BASE_MODE      : unsigned := to_unsigned(0,CLINKMODELEN);   -- 16 bit CLINK transfers
   constant CLINK_FULL_MODE      : unsigned := to_unsigned(1,CLINKMODELEN);   -- 64 bit CLINK transfers
   
   
   -- Pattern Generator Operational Mode Constants
   constant PG_STOP     : std_logic_vector(DIAGMODELEN-1 downto 0) := "0000";  -- Stop mode: forces a stop at the end of the next diag frame, triggering ignored
   constant PG_FRAME    : std_logic_vector(DIAGMODELEN-1 downto 0) := "0001";  -- Diagnostic mode: individual frame triggering mode
   constant PG_CAM_CNT  : std_logic_vector(DIAGMODELEN-1 downto 0) := "0010";  -- Diagnostic mode: Camera Frame simple pixel incrementation
   constant PG_CAM_VIS  : std_logic_vector(DIAGMODELEN-1 downto 0) := "0011";  -- Diagnostic mode: Camera Frame visible pattern
   constant PG_BSQ_XYZ  : std_logic_vector(DIAGMODELEN-1 downto 0) := "0100";  -- Diagnostic mode: BSQ DCube X,Y,Z counters
   constant PG_BIP_XYZ  : std_logic_vector(DIAGMODELEN-1 downto 0) := "0101";  -- Diagnostic mode: BIP DCube X,Y,Z counters
   constant PG_BIP_DIRAC: std_logic_vector(DIAGMODELEN-1 downto 0) := "0110";  -- Diagnostic mode: BIP DCube with Dirac for FFT tests (not yet implemented)
   constant PG_BSQ_COLD : std_logic_vector(DIAGMODELEN-1 downto 0) := "0111";  -- Diagnostic mode: BSQ DCube, cold BB
   constant PG_BSQ_HOT  : std_logic_vector(DIAGMODELEN-1 downto 0) := "1000";  -- Diagnostic mode: BSQ DCube, hot BB
   constant PG_BSQ_SCENE: std_logic_vector(DIAGMODELEN-1 downto 0) := "1001";  -- Diagnostic mode: BSQ DCube, real scene
   
   -- CLINK HEADER V4 Constants  (voir part 2 dans fichier excel)
   constant GEOPOS_LEN_V4          : integer := 104; -- nombre de bytes de la partie GEOPOSITIONNING dans le Header Clink v4 part2
   constant SPAREB_LEN_V4          : integer := 0; -- taille en bytes de SPARE_B dans le Header Clink v4 part2 
   
   constant NAV_DATA_REAL_V4_SIZE  : integer := GEOPOS_LEN_V4 - SPAREB_LEN_V4;
   
   constant SPAREA_LEN_V4          : integer := 32;   -- in bytes
   
   constant SPAREC_LEN_V4          : integer := 28;
   constant SPARED_LEN_V4          : integer := 28;
   constant SPAREE_LEN_V4          : integer := 32;
   constant SPAREF_LEN_V4          : integer := 56; 
   
   -- calcul
   constant SPAREAC_LEN_V4          : integer := SPAREA_LEN_V4 + SPAREC_LEN_V4;
   constant SPAREACD_LEN_V4         : integer := SPAREAC_LEN_V4 + SPARED_LEN_V4;
   constant SPAREACDE_LEN_V4        : integer := SPAREACD_LEN_V4 + SPAREE_LEN_V4;  
   constant SPAREACDEF_LEN_V4       : integer := SPAREACDE_LEN_V4 + SPAREF_LEN_V4;
   ------------------------------------------
   -- Types declarations
   ------------------------------------------
   
   type t_output_debug is
   record
      FPGA_ID : std_logic;
      Z : std_logic_vector(4 downto 0);
      Y : std_logic_vector(4 downto 0);
      X : std_logic_vector(4 downto 0);
   end record;
   
   type t_output_debug32 is
   record
      H : t_output_debug;
      L : t_output_debug;
   end record;
   
   type t_ddr_data21_debug is
   record
      P0 : std_logic_vector(20 downto 0);
      P1 : std_logic_vector(20 downto 0);
      P2 : std_logic_vector(20 downto 0);
      P3 : std_logic_vector(20 downto 0);
      P4 : std_logic_vector(20 downto 0);
      P5 : std_logic_vector(20 downto 0);
   end record;
   
   type t_RS232 is (CMD_40, CMD_41, CMD_42, CMD_43, CMD_44, CMD_50, CMD_60, CMD_61, CMD_62, CMD_92, CMD_93, CMD_94);
   
   type t_DIMM_CMD is (NOP, ACT, RD, WR, B_END, PRECH, RFRSH, LOAD, UNKNOWN);
   type DCUBE_HEADER_array is array (1 to DCUBE_HEADER_V2_size) of std_logic_vector(7 downto 0);   
   type DCUBE_HEADER_V2_array is array (1 to 12) of std_logic_vector(15 downto 0);
   type DCUBE_HEADER_V3_array is array (1 to DCUBE_HEADER_V3_size/2) of std_logic_vector(15 downto 0); -- new fixed part of header (external update)
   type DCUBE_FOOTER_V3_array is array (1 to DCUBE_FOOTER_V3_size/2) of std_logic_vector(15 downto 0); -- new status part of header (internal generation, may become footer)
   type DCUBE_FOOTER_V3_array8 is array (1 to DCUBE_FOOTER_V3_size) of std_logic_vector(7 downto 0); -- new status part of header (internal generation, may become footer)
   
   type ROIC_CLink_Header_array16 is array (1 to 18) of std_logic_vector(15 downto 0); -- This is the ROIC section in the CameraLink Header Part 2
   
   -- Version 4
   type DCUBE_Header_part1_array8_v4 is array (1 to DCUBE_part1_V4_size) of std_logic_vector(7 downto 0);
   type DCUBE_Header_part2_array8_v4 is array (1 to DCUBE_part2_V4_size) of std_logic_vector(7 downto 0);   
   
   type ROIC_CLink_Header_array16_v4 is array (1 to 32) of std_logic_vector(15 downto 0); -- This is the ROIC section in the CameraLink Header Part 2
   type DCUBE_Header_Part2_array_v4 is array (1 to DCUBE_part2_V4_size/2) of std_logic_vector(15 downto 0); -- new status part of header (internal generation, may become footer)
   type DCUBE_Header_Part1_array_v4 is array (1 to DCUBE_part1_V4_size/2) of std_logic_vector(15 downto 0);                                           
   type NAV_CLINK_Header_array16_v4 is array (1 to NAV_DATA_REAL_V4_SIZE/2) of std_logic_vector(15 downto 0); -- This is the NAV section in the CameraLink Header Part 2 (excluding SPARE_B
   
   type Camera_Link_Param_type is
   record
      LValSize    : unsigned(LVALLEN-1 downto 0);
      FValSize    : unsigned(FVALLEN-1 downto 0);
      HeaderSize  : unsigned(HEADERLEN-1 downto 0);
      LValPause   : unsigned(LPAUSELEN-1 downto 0);
      Clink_Mode  : std_logic_vector(CLINKMODELEN-1 downto 0);
   end record;
   
   type SpectralBand_Param_type is
   record
      Min   : unsigned(SBANDLEN-1 downto 0);
      Max   : unsigned(SBANDLEN-1 downto 0);
      Mode  : std_logic_vector(1 downto 0);
   end record;
   
   type VP30StatusInfo is
   record
      ExtTemp               : std_logic_vector(7 downto 0);
      IntTemp               : std_logic_vector(7 downto 0);
      Stat                  : std_logic_vector(31 downto 0);
   end record;
   
   type DPB_DCube_Header is -- These cubes are ALWAYS BIP, BSQ cubes start with ROIC_DCube_Header
   record
      DUI         : unsigned(DUILEN-1 downto 0); -- 4 bytes allocated for that field
      VP30Status  : VP30StatusInfo;    -- 8 bytes allocated for that field (for expansion)
      ROICHeader  : ROIC_DCube_Header; -- Info needed to populate the CameraLink Header
      ROICFooter  : ROIC_DCube_Footer; -- Info needed to populate the CameraLink Header
   end record;  
   
   type DPB_DCube_Header_v2_6 is -- These cubes are ALWAYS BIP, BSQ cubes start with ROIC_DCube_Header
   record
      DPBStatus         : std_logic_vector(DPBSTATLEN-1 downto 0);
      FirmwareVersion   : std_logic_vector(15 downto 0);
      FPGATemp          : std_logic_vector(7 downto 0);
      PCBTemp           : std_logic_vector(7 downto 0);
      PixelsReceivedCnt : unsigned(DUILEN-1 downto 0); -- 4 bytes allocated for that field      
      ROICHeader        : ROIC_DCube_Header_v2_6; -- Info needed to populate the CameraLink Header
      ROICFooter        : ROIC_DCube_Footer_v2_6; -- Info needed to populate the CameraLink Header
      NAVHeader         : NAV_DCube_Header_v2_6; -- Info needed to populate the CameraLink Header
   end record;
   constant DPB_DCube_Header_v2_6_32_LEN : natural := 5; -- Length including the header
   
   type DPB_DCube_Header_array16 is array (1 to 6 + ROIC_DCube_Header_array16'LENGTH + ROIC_DCube_Footer_array16'LENGTH) of std_logic_vector(15 downto 0);
   type DPB_DCube_Header_array32 is array (1 to 2 + ROIC_DCube_Header_array32'LENGTH + ROIC_DCube_Footer_array32'LENGTH) of std_logic_vector(31 downto 0);
   
   type DPB_DCube_Header_array32_v2_6 is array (1 to DPB_DCube_Header_v2_6_32_LEN + ROIC_DCube_Header_array32_v2_6'LENGTH + NAV_DCube_Header_array32_v2_6'LENGTH + ROIC_DCube_Footer_array32_v2_6'LENGTH) of std_logic_vector(31 downto 0);
   
   -- Pattern Generator Configuration
   type PatGenConfig is
   record
      DiagMode       : std_logic_vector(DIAGMODELEN-1 downto 0);  -- type of data frame to shoot.
      ZSize          : unsigned(ZLEN-1 downto 0);                 -- pixel count in z direction
      XSize          : unsigned(XLEN-1 downto 0);                 -- pixel count in x direction
      YSize          : unsigned(YLEN-1 downto 0);                 -- pixel count in y direction
      TagSize        : unsigned(TAGLEN-1 downto 0);               -- in BSQ data cube image mode (PG_BSQ_XYZ) number of pixels used by tag
      DiagSize       : unsigned(DIAGSIZELEN-1 downto 0);          -- number of succesive patterns to generate => 0= forever, 1-xxx = count
      PayloadSize    : unsigned(PLLEN-1 downto 0);                -- for filling frame ID header payload size value (24 bits)
      ImagePause     : unsigned(15 downto 0);                     -- Number of clock cycles to wait between each image, to trottle throughput.
      ROM_Z_START    : unsigned(15 downto 0);
      ROM_INIT_INDEX : unsigned(15 downto 0);
      IMGSIZE        : unsigned(IMGLEN-1 downto 0);
      
      Trig           : std_logic;                                 -- for triggering a pattern
      FrameType      : std_logic_vector(7 downto 0);              -- corresponds to frame ID header            
   end record;
   
   type patgen_array8 is array(1 to 34) of std_logic_vector(7 downto 0);   -- for RS232 transmition
   
   -- CameraLink board Configuration (from main controller)
   -- Note: Diagnostic mode settings are no longer appropriate in CLinkConfig.  However all array conversion
   -- functions support original array sizes so software needs no changes. The Mode and DiagSize fields
   -- are simply ignored
   type CLinkConfig is
   record
      Valid          : boolean; -- should pulse true for one clock after valid transmission to enable registering.
      -- CameraLink Settings
      LValSize       : unsigned(LVALLEN-1 downto 0);
      FValSize       : unsigned(FVALLEN-1 downto 0);
      HeaderSize     : unsigned(HEADERLEN-1 downto 0);
      LValPause      : unsigned(LPAUSELEN-1 downto 0);
      FramesPerCube  : unsigned(FRAMESPERCUBELEN-1 downto 0);
      CLinkMode      : unsigned(CLINKMODELEN-1 downto 0);
      HeaderVersion  : std_logic_vector(3 downto 0);
      -- Mode           : std_logic_vector(DIAGMODELEN-1 downto 0);  -- 0: Stop, 1: Normal, 2: Diagnostic #1, 3: Diagnostic #2
      -- DiagSize       : unsigned(DIAGSIZELEN-1 downto 0); -- range TBC
   end record;
   type CLinkConfig_array8 is array(1 to 38) of std_logic_vector(7 downto 0);   -- for RS232 transmition
   type CLinkConfig_array32 is array(1 to 10) of std_logic_vector(31 downto 0); -- for LocalLink transmition
   
   -- pragma translate_off
   -- DPConfig should only be used for simulation!
   type DPConfig is
   record
      ZSIZE       : unsigned(ZLEN-1 downto 0);
      XSIZE	      : unsigned(XLEN-1 downto 0);
      YSIZE		   : unsigned(YLEN-1 downto 0);
      IMGSIZE     : unsigned(IMGLEN-1 downto 0);
      TAGSIZE	   : unsigned(TAGLEN-1 downto 0);
      
      SB_Min      : unsigned(SBANDLEN-1 downto 0);
      SB_Max      : unsigned(SBANDLEN-1 downto 0);
      SB_Mode     : unsigned(1 downto 0);
      
      Interleave  : std_logic_vector(1 downto 0);
      Mode	      : std_logic_vector(DPMODELEN-1 downto 0);
      AVGSIZE	   : unsigned(AVGLEN-1 downto 0);
      DIAGSIZE    : unsigned(DIAGLEN-1 downto 0);
      
      BB_Temp     : unsigned(15 downto 0);
      Delta_OPD   : std_logic_vector(31 downto 0); -- float32 in fact
      Max_Temp    : unsigned(15 downto 0);
      --Gain_Exp    : signed(7 downto 0);
      --Off_Exp     : signed(7 downto 0); 
      SB_Min_Cal  : unsigned(SBANDLEN-1 downto 0);
      SB_Max_Cal  : unsigned(SBANDLEN-1 downto 0);      
   end record;
   -- pragma translate_on
   
   type DPConfig_array8 is array(1 to 70) of std_logic_vector(7 downto 0);
   type DPConfig_array32 is array(1 to 18) of std_logic_vector(31 downto 0);
   
   -- Data processing board Configuration (from main controller)
   type DPBConfig is
   record
      Camera_Link_Param    : Camera_Link_Param_type;
      SpectralBand_Param   : SpectralBand_Param_type;
      Datacube_Interleave  : std_logic_vector(1 downto 0);
      DP_Mode              : std_logic_vector(1 downto 0);
      Spare                : unsigned(7 downto 0);
      Fringe_Total         : unsigned(ZLEN-1 downto 0);
      XSIZE                : unsigned(XLEN-1 downto 0);
      YSIZE                : unsigned(YLEN-1 downto 0);
      IMGSIZE              : unsigned(IMGLEN-1 downto 0);
      TAGSIZE              : unsigned(TAGLEN-1 downto 0);
      AVGSIZE              : unsigned(AVGLEN-1 downto 0);
      HeaderVersion        : std_logic_vector(3 downto 0);
   end record;
   
   type VP7StatusInfo is
   record
      ExtTemp               : std_logic_vector(7 downto 0);
      IntTemp               : std_logic_vector(7 downto 0);
      Stat                  : std_logic_vector(31 downto 0);
   end record;
   
   -- Configuration for the module output_data_mem_read
   type MemReadConfigOld is
   record
      IMGSize           : unsigned(IMGLEN-1 downto 0);
      TAGSize           : unsigned(TAGLEN-1 downto 0);
      ZSize             : unsigned(ZLEN-1 downto 0);
      PAGE_SIZE         : unsigned(PAGELEN-1 downto 0);
      MemAdd            : std_logic_vector(AMAX downto 0); -- Only 256 Address Memory Zones
      MemInterleave     : std_logic_vector(1 downto 0);
      OutputInterleave  : std_logic_vector(1 downto 0);
      BitMode           : std_logic;
   end record;
   
   type MemReadConfig is
   record
      --IMGSIZE       : unsigned(IMGLEN-1 downto 0);
      ZSIZE         : unsigned(ZLEN-1 downto 0);
      PAGESIZE      : unsigned(PAGELEN-1 downto 0);
      PIXELNUM      : unsigned(IMGLEN-1 downto 0); -- Number of pixels to read
      INIT_ADD      : unsigned(AMAX downto 0);
      DDR_ADD_MAX   : unsigned(AMAX downto 0);
      CONTROL       : std_logic_vector(0 downto 0);
      CONFIG        : std_logic_vector(7 downto 0);
   end record;
   
   type MemWriteConfig is
   record
      IMGSIZE           : unsigned(IMGLEN-1 downto 0);
      IMGSIZE_M1        : unsigned(IMGLEN-1 downto 0);
      ZSIZE             : unsigned(ZLEN-1 downto 0);
      ZSIZE_M1          : unsigned(ZLEN-1 downto 0);
      ZSIZE_M1_D6_P1    : unsigned(ZLEN-3 downto 0);
      ZSIZE_M1_D8_P1    : unsigned(ZLEN-4 downto 0);
      LAST_PAGE_CNT_M1  : unsigned(2 downto 0); -- Number of valid images in the last ZBT page, minus 1.      
      TAGSIZE           : unsigned(TAGLEN-1 downto 0);
      AVGSIZE           : unsigned(AVGLEN-1 downto 0);
      INIT_ADD          : unsigned(AMAX downto 0);
      CONTROL           : std_logic_vector(0 downto 0);
      CONFIG            : std_logic_vector(7 downto 0);
   end record;
   
   type DiagConfig is
   record
      --Interleave     : std_logic_vector(1 downto 0);
      DP_Mode        : std_logic_vector(DPMODELEN-1 downto 0);
      ZSIZE          : unsigned(ZLEN-1 downto 0);
      XSIZE_ADJ      : unsigned(XLEN-1 downto 0);
      YSIZE          : unsigned(YLEN-1 downto 0);
      TAGSIZE        : unsigned(TAGLEN-1 downto 0);
      --AVGSIZE        : unsigned(AVGLEN-1 downto 0);
      DIAG_ACQ_NUM   : unsigned(9 downto 0);
      DATASIZE_M1    : unsigned(15 downto 0);
      ROM_Z_START    : unsigned(15 downto 0);
      ROM_INIT_INDEX : unsigned(15 downto 0);
      CONFIG         : std_logic_vector(7 downto 0);
   end record;
   
   type CalibConfig is
   record
      FRAMECNT       : unsigned(IMGLEN-1 downto 0) ; -- IMGSIZE without tags
      GAIN_EXPON     : std_logic_vector(7 downto 0);
      OFF_EXPON      : std_logic_vector(7 downto 0);
      EXTRA_EXPON    : std_logic_vector(7 downto 0);
      CONTROL        : std_logic_vector(1 downto 0);
      CONFIG         : std_logic_vector(1 downto 0);
      SB_Min         : unsigned(SBANDLEN-1 downto 0);
      SB_Max         : unsigned(SBANDLEN-1 downto 0);      
   end record;
   
   type DCUBE_FOOTER_V3 is
   record
      --Unused1                 : std_logic_vector(7 downto 0);
      DCA_SweepDirection      : std_logic;
      DCA_DataCubeID          : unsigned(22 downto 0);
      DCA_IntFramesCnt        : unsigned(31 downto 0);
      DCA_SampTrigsCnt        : unsigned(31 downto 0);
      DCA_ROICFirmwareVersion : std_logic_vector(15 downto 0);
      --SpareA                  : std_logic_vector(15 downto 0);
      DCA_ROICStatus          : std_logic_vector(15 downto 0);
      DCA_FOVStartX           : unsigned(15 downto 0);
      DCA_FOVStartY           : unsigned(15 downto 0);
      DCA_ZPDPosition         : unsigned(31 downto 0);
      DCA_MaxFPACount         : unsigned(15 downto 0);
      DCA_TimeStamp           : unsigned(31 downto 0);
      --SpareB                  : std_logic_vector(31 downto 0);
      --Unused2                 : std_logic_vector(7 downto 0);
      DCA_FPGA1_Status        : VP30StatusInfo;
      --SpareC                  : std_logic_vector(31 downto 0);
      --Unused3                 : std_logic_vector(7 downto 0);
      DCA_FPGA2_Status        : VP30StatusInfo;
      --SpareD                  : std_logic_vector(31 downto 0);
      --Unused4                 : std_logic_vector(7 downto 0);
      DCA_FPGA3_Status        : VP7StatusInfo;
      DCA_DUI                 : unsigned(31 downto 0);
      DCA_DPBFirmwareVersion  : std_logic_vector(15 downto 0);
      --SpareE                  : std_logic_vector(159 downto 0);
   end record;
   
   --   type DCUBE_Header_Part2_v4 is
   --   record
   --      --Unused1                 : std_logic_vector(7 downto 0);
   --      DCA_SweepDirection      : std_logic;
   --      DCA_DataCubeID          : unsigned(22 downto 0);
   --      DCA_IntFramesCnt        : unsigned(31 downto 0);
   --      DCA_SampTrigsCnt        : unsigned(31 downto 0);
   --      DCA_ROICFirmwareVersion : std_logic_vector(15 downto 0);
   --      --SpareA                  : std_logic_vector(15 downto 0);
   --      DCA_ROICStatus          : std_logic_vector(15 downto 0);
   --      DCA_FOVStartX           : unsigned(15 downto 0);
   --      DCA_FOVStartY           : unsigned(15 downto 0);
   --      DCA_ZPDPosition         : unsigned(31 downto 0);
   --      DCA_MaxFPACount         : unsigned(15 downto 0);
   --      DCA_TimeStamp           : unsigned(31 downto 0);
   --      --SpareB                  : std_logic_vector(31 downto 0);
   --      --Unused2                 : std_logic_vector(7 downto 0);
   --      DCA_FPGA1_Status        : VP30StatusInfo;
   --      --SpareC                  : std_logic_vector(31 downto 0);
   --      --Unused3                 : std_logic_vector(7 downto 0);
   --      DCA_FPGA2_Status        : VP30StatusInfo;
   --      --SpareD                  : std_logic_vector(31 downto 0);
   --      --Unused4                 : std_logic_vector(7 downto 0);
   --      DCA_FPGA3_Status        : VP7StatusInfo;
   --      DCA_DUI                 : unsigned(31 downto 0);
   --      DCA_DPBFirmwareVersion  : std_logic_vector(15 downto 0);
   --      --SpareE                  : std_logic_vector(159 downto 0);
   --   end record;
   
   
   ------------------------------------------
   -- Project constants
   ------------------------------------------
   constant RIO_latency : integer := 80;
   constant MODE_delay  : integer := 100;
   
   constant DPBConfig_size : integer := DPBConfig_array'LENGTH;
   
   --   constant VP30StatusInfo_default : VP30StatusInfo :=
   --   (x"00", x"00", DPB_VERSION & x"000000");
   
   constant VP7StatusInfo_default : VP7StatusInfo :=
   (x"00", x"00", CLINK_VERSION & x"000000");
   
   constant DCUBE_HEADER_array_default : DCUBE_HEADER_array :=
   (X"00", X"01", X"02", X"03", X"04", X"05", X"06", X"07", X"08", X"09", X"0A", X"0B", X"0C", X"0D", X"0E", X"0F",
   X"10", X"11", X"12", X"13", X"14", X"15", X"16", X"17", X"18", X"19", X"1A", X"1B", X"1C", X"1D", X"1E", X"1F",
   X"20", X"21", X"22", X"23", X"24", X"25", X"26", X"27", X"28", X"29", X"2A", X"2B", X"2C", X"2D", X"2E", X"2F",
   X"30", X"31", X"32", X"33", X"34", X"35", X"36", X"37", X"38", X"39", X"3A", X"3B", X"3C", X"3D", X"3E", X"3F",
   X"40", X"41", X"42", X"43", X"44", X"45", X"46", X"47", X"48", X"49", X"4A", X"4B", X"4C", X"4D", X"4E", X"4F",
   X"50", X"51", X"52", X"53", X"54", X"55", X"56", X"57", X"58", X"59", X"5A", X"5B", X"5C", X"5D", X"5E", X"5F",
   X"60", X"61", X"62", X"63", X"64", X"65", X"66", X"67", X"68", X"69", X"6A", X"6B", X"6C", X"6D", X"6E", X"6F",
   X"70", X"71", X"72", X"73", X"74", X"75", X"76", X"77", X"78", X"79", X"7A", X"7B", X"7C", X"7D", X"7E", X"7F",
   X"80", X"81", X"82", X"83", X"84", X"85", X"86", X"87", X"88", X"89", X"8A", X"8B", X"8C", X"8D", X"8E", X"8F",
   X"90", X"91", X"92", X"93", X"94", X"95", X"96", X"97", X"98", X"99", X"9A", X"9B", X"9C", X"9D", X"9E", X"9F",
   X"A0", X"A1", X"A2", X"A3", X"A4", X"A5", X"A6", X"A7", X"A8", X"A9", X"AA", X"AB", X"AC", X"AD", X"AE", X"AF",
   X"B0", X"B1", X"B2", X"B3", X"B4", X"B5", X"B6", X"B7", X"B8", X"B9", X"BA", X"BB", X"BC", X"BD", X"BE", X"BF",
   X"C0", X"C1", X"C2", X"C3", X"C4", X"C5", X"C6", X"C7", X"C8", X"C9", X"CA", X"CB", X"CC", X"CD", X"CE", X"CF",
   X"D0", X"D1", X"D2", X"D3", X"D4", X"D5", X"D6", X"D7", X"D8", X"D9", X"DA", X"DB", X"DC", X"DD", X"DE", X"DF",
   X"E0", X"E1", X"E2", X"E3", X"E4", X"E5", X"E6", X"E7", X"E8", X"E9", X"EA", X"EB", X"EC", X"ED", X"EE", X"EF",
   X"F0", X"F1", X"F2", X"F3", X"F4", X"F5", X"F6", X"F7", X"F8", X"F9", X"FA", X"FB", X"FC", X"FD", X"FE", X"FF",
   X"00", X"01", X"02", X"03", X"04", X"05", X"06", X"07", X"08", X"09", X"0A", X"0B", X"0C", X"0D", X"0E", X"0F",
   X"10", X"11", X"12", X"13", X"14", X"15", X"16", X"17", X"18", X"19", X"1A", X"1B", X"1C", X"1D", X"1E", X"1F",
   X"20", X"21", X"22", X"23", X"24", X"25", X"26", X"27", X"28", X"29", X"2A", X"2B", X"2C", X"2D", X"2E", X"2F",
   X"30", X"31", X"32", X"33", X"34", X"35", X"36", X"37", X"38", X"39", X"3A", X"3B", X"3C", X"3D", X"3E", X"3F",
   X"40", X"41", X"42", X"43", X"44", X"45", X"46", X"47", X"48", X"49", X"4A", X"4B", X"4C", X"4D", X"4E", X"4F",
   X"50", X"51", X"52", X"53", X"54", X"55", X"56", X"57", X"58", X"59", X"5A", X"5B", X"5C", X"5D", X"5E", X"5F",
   X"60", X"61", X"62", X"63", X"64", X"65", X"66", X"67", X"68", X"69", X"6A", X"6B", X"6C", X"6D", X"6E", X"6F",
   X"70", X"71", X"72", X"73", X"74", X"75", X"76", X"77", X"78", X"79", X"7A", X"7B", X"7C", X"7D", X"7E", X"7F",
   X"80", X"81", X"82", X"83", X"84", X"85", X"86", X"87", X"88", X"89", X"8A", X"8B", X"8C", X"8D", X"8E", X"8F",
   X"90", X"91", X"92", X"93", X"94", X"95", X"96", X"97", X"98", X"99", X"9A", X"9B", X"9C", X"9D", X"9E", X"9F",
   X"A0", X"A1", X"A2", X"A3", X"A4", X"A5", X"A6", X"A7", X"A8", X"A9", X"AA", X"AB", X"AC", X"AD", X"AE", X"AF",
   X"B0", X"B1", X"B2", X"B3", X"B4", X"B5", X"B6", X"B7", X"B8", X"B9", X"BA", X"BB", X"BC", X"BD", X"BE", X"BF",
   X"C0", X"C1", X"C2", X"C3", X"C4", X"C5", X"C6", X"C7", X"C8", X"C9", X"CA", X"CB", X"CC", X"CD", X"CE", X"CF",
   X"D0", X"D1", X"D2", X"D3", X"D4", X"D5", X"D6", X"D7", X"D8", X"D9", X"DA", X"DB", X"DC", X"DD", X"DE", X"DF",
   X"E0", X"E1", X"E2", X"E3", X"E4", X"E5", X"E6", X"E7", X"E8", X"E9", X"EA", X"EB", X"EC", X"ED", X"EE", X"EF",
   X"F0", X"F1", X"F2", X"F3", X"F4", X"F5", X"F6", X"F7", X"F8", X"F9", X"FA", X"FB", X"FC", X"FD", X"FE", X"FF");
   constant DCUBE_HEADER_V3_array_default : DCUBE_HEADER_V3_array :=
   (X"0001", X"0203", X"0405", X"0607", X"0809", X"0A0B", X"0C0D", X"0E0F",
   X"1011", X"1213", X"1415", X"1617", X"1819", X"1A1B", X"1C1D", X"1E1F",
   X"2021", X"2223", X"2425", X"2627", X"2829", X"2A2B", X"2C2D", X"2E2F",
   X"3031", X"3233", X"3435", X"3637", X"3839", X"3A3B", X"3C3D", X"3E3F",
   X"4041", X"4243", X"4445", X"4647", X"4849", X"4A4B", X"4C4D", X"4E4F",
   X"5051", X"5253", X"5455", X"5657", X"5859", X"5A5B", X"5C5D", X"5E5F",
   X"6061", X"6263", X"6465", X"6667", X"6869", X"6A6B", X"6C6D", X"6E6F",
   X"7071", X"7273", X"7475", X"7677", X"7879", X"7A7B", X"7C7D", X"7E7F",
   X"8081", X"8283", X"8485", X"8687", X"8889", X"8A8B", X"8C8D", X"8E8F",
   X"9091", X"9293", X"9495", X"9697", X"9899", X"9A9B", X"9C9D", X"9E9F",
   X"A0A1", X"A2A3", X"A4A5", X"A6A7", X"A8A9", X"AAAB", X"ACAD", X"AEAF",
   X"B0B1", X"B2B3", X"B4B5", X"B6B7", X"B8B9", X"BABB", X"BCBD", X"BEBF",
   X"C0C1", X"C2C3", X"C4C5", X"C6C7", X"C8C9", X"CACB", X"CCCD", X"CECF",
   X"D0D1", X"D2D3", X"D4D5", X"D6D7", X"D8D9", X"DADB", X"DCDD", X"DEDF",
   X"E0E1", X"E2E3", X"E4E5", X"E6E7", X"E8E9", X"EAEB", X"ECED", X"EEEF",
   X"F0F1", X"F2F3", X"F4F5", X"F6F7", X"F8F9", X"FAFB", X"FCFD", X"FEFF",
   X"0001", X"0203", X"0405", X"0607", X"0809", X"0A0B", X"0C0D", X"0E0F",
   X"1011", X"1213", X"1415", X"1617", X"1819", X"1A1B", X"1C1D", X"1E1F",
   X"2021", X"2223", X"2425", X"2627", X"2829", X"2A2B", X"2C2D", X"2E2F",
   X"3031", X"3233", X"3435", X"3637", X"3839", X"3A3B", X"3C3D", X"3E3F",
   X"4041", X"4243", X"4445", X"4647", X"4849", X"4A4B", X"4C4D", X"4E4F",
   X"5051", X"5253", X"5455", X"5657", X"5859", X"5A5B", X"5C5D", X"5E5F",
   X"6061", X"6263", X"6465", X"6667", X"6869", X"6A6B", X"6C6D", X"6E6F",
   X"7071", X"7273", X"7475", X"7677", X"7879", X"7A7B", X"7C7D", X"7E7F",
   X"8081", X"8283", X"8485", X"8687", X"8889", X"8A8B", X"8C8D", X"8E8F",
   X"9091", X"9293", X"9495", X"9697", X"9899", X"9A9B", X"9C9D", X"9E9F",
   X"A0A1", X"A2A3", X"A4A5", X"A6A7", X"A8A9", X"AAAB", X"ACAD", X"AEAF",
   X"B0B1", X"B2B3", X"B4B5", X"B6B7", X"B8B9", X"BABB", X"BCBD", X"BEBF",
   X"C0C1", X"C2C3", X"C4C5", X"C6C7", X"C8C9", X"CACB", X"CCCD", X"CECF",
   X"D0D1", X"D2D3", X"D4D5", X"D6D7", X"D8D9", X"DADB", X"DCDD", X"DEDF",
   X"E0E1", X"E2E3", X"E4E5", X"E6E7", X"E8E9", X"EAEB", X"ECED", X"EEEF",
   X"F0F1", X"F2F3", X"F4F5", X"F6F7", X"F8F9", X"FAFB", X"FCFD", X"FEFF");
   
   constant DCUBE_FOOTER_V3_array_default : DCUBE_FOOTER_V3_array :=
   (X"0001", X"0203", X"0405", X"0607", X"0809", X"0A0B", X"0C0D", X"0E0F",
   X"1011", X"1213", X"1415", X"1617", X"1819", X"1A1B", X"1C1D", X"1E1F",
   X"2021", X"2223", X"2425", X"2627", X"2829", X"2A2B", X"2C2D", X"2E2F",
   X"3031", X"3233", X"3435", X"3637", X"3839", X"3A3B", X"3C3D", X"3E3F",
   X"4041", X"4243", X"4445", X"4647", X"4849", X"4A4B", X"4C4D", X"4E4F",
   X"5051", X"5253", X"5455", X"5657");
   ------------------------------------------
   -- *** FUNCTIONS DECLARATIONS***
   ------------------------------------------
   function to_DPBConfig_array (a: DPBConfig) return DPBConfig_array;
   --function to_DPBConfig (a: DPBConfig_array; FPGA_ID: std_logic) return DPBConfig;
   
   -- pragma translate_off
   function to_DPBConfig (a: DPConfig; b: CLinkConfig) return DPBConfig;
   function to_CLinkConfig_array8 (a: CLinkConfig) return CLinkConfig_array8;
   -- pragma translate_on
   
   function to_CLinkConfig (a: CLinkConfig_array8; ValidConfig: boolean) return CLinkConfig;
   function to_CLinkConfig_array32 (a: CLinkConfig) return CLinkConfig_array32;
   function to_CLinkConfig (a: CLinkConfig_array32; ValidConfig: boolean) return CLinkConfig;
   function to_CLinkConfig (a: DPBConfig) return CLinkConfig;   -- For backward testbench compatibility
   
   -- pragma translate_off
   function to_DPConfig_array8 (a: DPConfig) return DPConfig_array8;
   function to_DPConfig_array8 (a: DPConfig; MissingImages : integer) return DPConfig_array8;
   function to_DPConfig (a: DPConfig_array8) return DPConfig;   
   function to_DPConfig_array32 (a: DPConfig) return DPConfig_array32;
   function to_DPConfig_array32 (a: DPConfig; MissingImages : integer) return DPConfig_array32;
   function to_DPConfig (a: DPBConfig; Mode : std_logic_vector) return DPConfig;   -- For backward testbench compatibility
   function to_DCUBE_HEADER_array (a: DPConfig; b: CLinkConfig) return DCUBE_HEADER_array;
   function to_DCUBE_Header_part1_array8_v4(a: DPConfig; b: CLinkConfig; SamplingPeriodNumerator: std_logic_vector) return DCUBE_Header_part1_array8_v4;
   function to_output_debug(a: std_logic_vector(15 downto 0)) return t_output_debug;
   function to_output_debug32(a: std_logic_vector(31 downto 0)) return t_output_debug32;
   function to_ddr_data21_debug(a: std_logic_vector(127 downto 0)) return t_ddr_data21_debug;
   -- pragma translate_on
   
   function to_ROIC_CLink_Header_array16(h: ROIC_DCube_Header; f: ROIC_DCube_Footer) return ROIC_CLink_Header_array16;
   function to_ROIC_CLink_Header_array16(h: ROIC_DCube_Header) return ROIC_CLink_Header_array16;
   function to_DCUBE_FOOTER_V3_array (a, b : DPB_DCube_Header; c : VP7StatusInfo) return DCUBE_FOOTER_V3_array;
   function to_DCUBE_FOOTER_V3_array (a: ROIC_DCube_Header; c : VP7StatusInfo) return DCUBE_FOOTER_V3_array;
   -- CLINK_header v4
   function to_DCUBE_Header_Part2_array_V4 (a, b : DPB_DCube_Header_v2_6; c : VP7StatusInfo; DP_Present: std_logic) return DCUBE_Header_Part2_array_V4;
   function to_ROIC_CLink_Header_array16_v4(h: ROIC_DCube_Header_v2_6;f: ROIC_DCube_Footer_v2_6; DP_Present :std_logic) return ROIC_CLink_Header_array16_v4;
   --function to_DCUBE_part2_V4_array (a: ROIC_DCube_Header_v2_6; c : VP7StatusInfo) return DCUBE_part2_V4_array;
   -- overloaded functions to standardize calling of similar things
   function to_std_logic_vector (a: VP7StatusInfo) return std_logic_vector;
   function to_std_logic_vector (a: VP30StatusInfo) return std_logic_vector;
   function to_VP30StatusInfo (a: std_logic_vector) return VP30StatusInfo;
   function to_VP7StatusInfo (a: std_logic_vector) return VP7StatusInfo;
   function status_latch (new_status,old_status: VP30StatusInfo) return VP30StatusInfo;
   function status_latch (new_status,old_status: VP7StatusInfo) return VP7StatusInfo;
   function to_DCUBE_FOOTER_V3 (b: DCUBE_FOOTER_V3_array) return DCUBE_FOOTER_V3;
   --function to_DCUBE_Header_Part2_v4 (b: DCUBE_Header_Part2_array_v4) return DCUBE_Header_Part2_v4;
   function to_DPB_DCube_Header(a: unsigned(DUILEN-1 downto 0); b: VP30StatusInfo; c: ROIC_DCube_Header; d: ROIC_DCube_Footer) return DPB_DCube_Header;
   function to_DPB_DCube_Header(a: DPB_DCube_Header_array16) return DPB_DCube_Header;
   
   function to_DPB_DCube_Header(a: DPB_DCube_Header_array32) return DPB_DCube_Header;
   function to_DPB_DCube_Header_array32(a: DPB_DCube_Header) return DPB_DCube_Header_array32; 
   
   function to_DPB_DCube_Header_v2_6(a: DPB_DCube_Header_array32_v2_6) return DPB_DCube_Header_v2_6;
   function to_DPB_DCube_Header_array32_v2_6(a: DPB_DCube_Header_v2_6) return DPB_DCube_Header_array32_v2_6;
   
   function to_PatGenConfig (a: patgen_array8; ValidConfig: boolean) return PatGenConfig;
   -- pragma translate_off
   function to_patgen_array8 (a: PatGenConfig) return patgen_array8;
   -- pragma translate_on
   function to_NAV_CLINK_Header_array16_v4(h: NAV_DCube_Header_v2_6) return NAV_CLINK_Header_array16_v4;
   
end DPB_Define;

------------------------------------------
-- *** ADMET_DEFINE PACKAGE BODY***
------------------------------------------
package body DPB_Define is
   
   function to_DPBConfig_array (a: DPBConfig) return DPBConfig_array is
      variable y: DPBConfig_array;
   begin
      y(1) := X"00";
      y(2) := X"00";
      y(3) := std_logic_vector(a.Camera_Link_Param.LValSize(15 downto 8));
      y(4) := std_logic_vector(a.Camera_Link_Param.LValSize(7 downto 0));
      y(5) := X"00";
      y(6) := X"00";
      y(7) := std_logic_vector(a.Camera_Link_Param.FValSize(15 downto 8));
      y(8) := std_logic_vector(a.Camera_Link_Param.FValSize(7 downto 0));
      y(9)  := std_logic_vector(a.Camera_Link_Param.HeaderSize(15 downto 8));
      y(10) := std_logic_vector(a.Camera_Link_Param.HeaderSize(7 downto 0));
      y(11) := std_logic_vector(a.Camera_Link_Param.LValPause(15 downto 8));
      y(12) := std_logic_vector(a.Camera_Link_Param.LValPause(7 downto 0));
      y(13) := std_logic_vector(a.SpectralBand_Param.Min(15 downto 8));
      y(14) := std_logic_vector(a.SpectralBand_Param.Min(7 downto 0));
      y(15) := std_logic_vector(a.TAGSIZE);
      y(16) := "00" & std_logic_vector(a.AVGSIZE);
      y(17) := std_logic_vector(a.SpectralBand_Param.Max(15 downto 8));
      y(18) := std_logic_vector(a.SpectralBand_Param.Max(7 downto 0));
      y(19) := "00" & a.HeaderVersion & a.SpectralBand_Param.Mode;
      y(20) := "000000" & a.Datacube_Interleave;
      y(21) := "000000" & a.DP_Mode;
      y(22) := std_logic_vector(a.Spare);
      y(23) := std_logic_vector(a.Fringe_Total(23 downto 16));
      y(24) := std_logic_vector(a.Fringe_Total(15 downto 8));
      y(25) := std_logic_vector(a.Fringe_Total(7 downto 0));
      y(26) := "000000" & std_logic_vector(a.XSIZE(9 downto 8));
      y(27) := std_logic_vector(a.XSIZE(7 downto 0));
      y(28) := "000000" & std_logic_vector(a.YSIZE(9 downto 8));
      y(29) := std_logic_vector(a.YSIZE(7 downto 0));
      return y;
   end to_DPBConfig_array;
   
   --   function to_DPBConfig (a: DPBConfig_array; FPGA_ID: std_logic) return DPBConfig is
   --      variable y: DPBConfig;
   --      variable XSIZE_adjust : integer range 0 to 1;
   --   begin
   --      y.Camera_Link_Param.LValSize := unsigned(a(3)) & unsigned(a(4));
   --      y.Camera_Link_Param.FValSize := unsigned(a(7)) & unsigned(a(8));
   --      y.Camera_Link_Param.HeaderSize := unsigned(a(9)) & unsigned(a(10));
   --      y.Camera_Link_Param.LValPause := unsigned(a(11)) & unsigned(a(12));
   --      y.SpectralBand_Param.Min := unsigned(a(13)) & unsigned(a(14));
   --      y.TAGSIZE := unsigned(a(15));
   --      y.AVGSIZE := unsigned(a(16)(5 downto 0));
   --      y.SpectralBand_Param.Max := unsigned(a(17)) & unsigned(a(18));
   --      y.HeaderVersion := a(19)(5 downto 2);
   --      y.SpectralBand_Param.Mode := a(19)(1 downto 0);
   --      y.Datacube_Interleave := a(20)(1 downto 0);
   --      y.DP_Mode := a(21)(y.DP_Mode'LENGTH-1 downto 0);
   --      y.Spare := unsigned(a(22));
   --      y.Fringe_Total := unsigned(a(23)) & unsigned(a(24)) & unsigned(a(25));
   --      y.XSIZE := unsigned(a(26)(1 downto 0)) & unsigned(a(27));
   --      y.YSIZE := unsigned(a(28)(1 downto 0)) & unsigned(a(29));
   --      if FPGA_ID = '0' then
   --         XSIZE_adjust := 1;
   --      else
   --         XSIZE_adjust := 0;
   --      end if;
   --      y.IMGSIZE := resize(((y.XSIZE+XSIZE_adjust)/2) * y.YSIZE, y.IMGSIZE'LENGTH);
   --      if y.AVGSIZE = 0 then
   --         y.AVGSIZE := to_unsigned(1, y.AVGSIZE'LENGTH);
   --      end if;
   --      return y;
   --   end to_DPBConfig;
   
   -- pragma translate_off
   function to_DPBConfig (a: DPConfig; b: CLinkConfig) return DPBConfig is
      variable y: DPBConfig;
   begin
      y.Datacube_Interleave := a.Interleave;
      y.DP_Mode := "00";
      y.XSIZE := a.XSIZE;
      y.YSIZE := a.YSIZE;
      y.Fringe_Total := a.ZSIZE;
      y.IMGSIZE := a.IMGSIZE;
      y.TAGSIZE := a.TAGSIZE;
      y.AVGSIZE := a.AVGSIZE;
      y.SpectralBand_Param.Mode := std_logic_vector(a.SB_Mode);
      y.SpectralBand_Param.Min := a.SB_Min;
      y.SpectralBand_Param.Max := a.SB_Max;
      y.Camera_Link_Param.LValSize :=   b.LValSize;
      y.Camera_Link_Param.FValSize :=   b.FValSize;
      y.Camera_Link_Param.HeaderSize := b.HeaderSize;
      y.Camera_Link_Param.LValPause :=  b.LValPause;
      return y;
      
   end to_DPBConfig;
   -- pragma translate_on
   
   -- translate_off
   function to_CLinkConfig_array8 (a: CLinkConfig) return CLinkConfig_array8 is
      variable y : CLinkConfig_array8;
      variable data32 : unsigned(31 downto 0);
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 9; -- In 32-bit elements
      constant PayloadSizeInBytes : integer := PayloadSize*4;
   begin
      y(1) := x"60";
      y(2) := std_logic_vector(to_unsigned(PayloadSizeInBytes,8)); -- Payload size
      
      for i in 1 to PayloadSize loop
         case i is
            when 1 => data32 := resize(a.LValSize, 32);
            when 2 => data32 := resize(a.FValSize, 32);
            when 3 => data32 := resize(a.HeaderSize, 32);
            when 4 => data32 := resize(a.LValPause, 32);
            when 5 => data32 := resize(a.FramesPerCube, 32);
            when 6 => data32 := resize(unsigned(a.CLinkMode), 32);
            when 7 => data32 := resize(unsigned(a.HeaderVersion), 32);
            when 8 => data32 := (others => '0');
            when 9 => data32 := (others => '0');
            -- when 8 => data32 := resize(unsigned(a.Mode), 32);
            -- when 9 => data32 := resize(a.DiagSize, 32);
         end case;
         data32_slv := std_logic_vector(data32);
         y(i*4-3 + 2) := data32_slv(31 downto 24); -- MSB
         y(i*4-2 + 2) := data32_slv(23 downto 16);
         y(i*4-1 + 2) := data32_slv(15 downto 8);
         y(i*4 + 2)   := data32_slv(7 downto 0);-- LSB
      end loop;
      
      return y;
   end to_CLinkConfig_array8;
   -- translate_on
   
   function to_CLinkConfig (a: CLinkConfig_array8; ValidConfig: boolean) return CLinkConfig is
      variable y : CLinkConfig;
      variable data32 : unsigned(31 downto 0);
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 9;
   begin
      -- pragma translate_off
      assert a(1) = x"60" report "Wrong header received, expected 0x60" severity ERROR;
      if ValidConfig then
         assert (to_integer(unsigned(a(2))) = CLinkConfig_array8'LENGTH-2) report "Wrong payload size received for command 0x60" severity ERROR;
      end if;
      -- pragma translate_on
      
      for i in 1 to PayloadSize loop
         data32_slv := a(i*4-3 + 2) & a(i*4-2 + 2) & a(i*4-1 + 2) & a(i*4 + 2);
         data32 := unsigned(data32_slv);
         
         case i is
            when 1 => y.LValSize       := resize(data32, LVALLEN);
            when 2 => y.FValSize       := resize(data32, FVALLEN);
            when 3 => y.HeaderSize     := resize(data32, HEADERLEN);
            when 4 => y.LValPause      := resize(data32, LPAUSELEN);
            when 5 => y.FramesPerCube  := resize(data32, FRAMESPERCUBELEN);
            when 6 => y.CLinkMode      := resize(data32, CLINKMODELEN);
            when 7 => y.HeaderVersion  := std_logic_vector(resize(data32, y.HeaderVersion'LENGTH));
            when 8 => null;
            when 9 => null;
            -- when 8 => y.Mode           := std_logic_vector(resize(data32, y.Mode'LENGTH         ));
            -- when 9 => y.DiagSize       := resize(data32, y.DiagSize'LENGTH);
         end case;
      end loop;
      
      y.Valid := ValidConfig;
      
      return y;
   end to_CLinkConfig;
   
   function to_CLinkConfig_array32 (a: CLinkConfig) return CLinkConfig_array32 is
      variable y : CLinkConfig_array32;
      constant PayloadSize : integer := 9; -- In 32-bit elements
   begin
      y(1) := x"60" & std_logic_vector(to_unsigned(PayloadSize,24)); -- Payload size
      y(2) := std_logic_vector(resize(a.LValSize, 32));
      y(3) := std_logic_vector(resize(a.FValSize, 32));
      y(4) := std_logic_vector(resize(a.HeaderSize, 32));
      y(5) := std_logic_vector(resize(a.LValPause, 32));
      y(6) := std_logic_vector(resize(a.FramesPerCube, 32));
      y(7) := std_logic_vector(resize(unsigned(a.CLinkMode), 32));
      y(8) := std_logic_vector(resize(unsigned(a.HeaderVersion), 32));
      -- y(9) := std_logic_vector(resize(unsigned(a.Mode), 32));
      -- y(10):= std_logic_vector(resize(a.DiagSize, 32));
      return y;
   end to_CLinkConfig_array32;
   
   function to_CLinkConfig (a: CLinkConfig_array32; ValidConfig: boolean) return CLinkConfig is
      variable y : CLinkConfig;
      constant PayloadSize : integer := 9;
   begin
      -- pragma translate_off
      assert a(1)(31 downto 24) = x"60" report "Wrong header received, expected 0x60" severity ERROR;
      if ValidConfig then
         assert (to_integer(unsigned(a(1)(23 downto 0))) = CLinkConfig_array32'LENGTH-1) report "Wrong payload size received for command 0x60" severity ERROR;
      end if;
      -- pragma translate_on
      
      y.LValSize       := resize(unsigned(a(2)), LVALLEN);
      y.FValSize       := resize(unsigned(a(3)), FVALLEN);
      y.HeaderSize     := resize(unsigned(a(4)), HEADERLEN);
      y.LValPause      := resize(unsigned(a(5)), LPAUSELEN);
      y.FramesPerCube  := resize(unsigned(a(6)), FRAMESPERCUBELEN);
      y.CLinkMode      := resize(unsigned(a(7)), CLINKMODELEN);
      y.HeaderVersion  := std_logic_vector(resize(unsigned(a(8)), y.HeaderVersion'LENGTH));
      -- y.Mode           := std_logic_vector(resize(unsigned(a(9)), y.Mode'LENGTH));
      -- y.DiagSize       := resize(unsigned(a(10)), y.DiagSize'LENGTH);
      y.Valid          := ValidConfig;
      
      return y;
   end to_CLinkConfig;
   
   
   function to_CLinkConfig (a: DPBConfig) return CLinkConfig is
      variable y : CLinkConfig;
   begin
      y.LValSize       := a.Camera_Link_Param.LValSize;
      y.FValSize       := a.Camera_Link_Param.FValSize;
      y.HeaderSize     := a.Camera_Link_Param.HeaderSize;
      y.LValPause      := a.Camera_Link_Param.LValPause;
      y.FramesPerCube  := x"0001"; -- No multi frames
      y.CLinkMode      := (others => '0');
      y.HeaderVersion  := x"3";
      -- y.Mode           := "001"; -- Normal mode
      -- y.DiagSize       := x"0001";
      return y;
   end to_CLinkConfig;
   
   -- pragma translate_off
   function to_DPConfig_array8 (a: DPConfig) return DPConfig_array8 is
      variable y : DPConfig_array8;
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 17; -- In 32-bit elements
      constant PayloadSizeInBytes : integer := PayloadSize*4;
   begin
      y(1) := x"61";
      y(2) := std_logic_vector(to_unsigned(PayloadSizeInBytes,8)); -- Payload size
      
      for i in 1 to PayloadSize loop
         case i is
            when 1  => data32_slv := std_logic_vector(resize(a.ZSIZE	   , 32));
            when 2  => data32_slv := std_logic_vector(resize(a.XSIZE	   , 32));
            when 3  => data32_slv := std_logic_vector(resize(a.YSIZE		, 32));
            when 4  => data32_slv := std_logic_vector(resize(a.IMGSIZE  , 32));
            when 5  => data32_slv := std_logic_vector(resize(a.TAGSIZE	, 32));
            when 6  => data32_slv := std_logic_vector(resize(a.SB_Min   , 32));
            when 7  => data32_slv := std_logic_vector(resize(a.SB_Max   , 32));
            when 8  => data32_slv := std_logic_vector(resize(a.SB_Mode  , 32));
            when 9  => data32_slv := std_logic_vector(resize(unsigned(a.Interleave) , 32));
            when 10 => data32_slv := std_logic_vector(resize(unsigned(a.Mode)       , 32));
            when 11 => data32_slv := std_logic_vector(resize(a.AVGSIZE	  , 32));
            when 12 => data32_slv := std_logic_vector(resize(a.DIAGSIZE   , 32));
            when 13 => data32_slv := std_logic_vector(resize(a.BB_Temp    , 32));
            when 14 => data32_slv := std_logic_vector(resize(unsigned(a.Delta_OPD)  , 32));
            when 15 => data32_slv := std_logic_vector(resize(a.Max_Temp   , 32));
            when 16 => data32_slv := std_logic_vector(resize(a.SB_Min_Cal   , 32));
            when 17 => data32_slv := std_logic_vector(resize(a.SB_Max_Cal    , 32));
            --when 18 => data32_slv := std_logic_vector(resize(a.Lh_Exp     , 32));
            --when 19 => data32_slv := std_logic_vector(resize(a.DLbb_Exp   , 32));
         end case;
         
         y(i*4-3 + 2) := data32_slv(31 downto 24); -- MSB
         y(i*4-2 + 2) := data32_slv(23 downto 16);
         y(i*4-1 + 2) := data32_slv(15 downto 8);
         y(i*4 + 2)   := data32_slv(7 downto 0);-- LSB
      end loop;
      
      return y;
   end to_DPConfig_array8;  
   
   function to_DPConfig_array8 (a: DPConfig; MissingImages : integer) return DPConfig_array8 is
      variable y : DPConfig_array8;
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 17; -- In 32-bit elements
      constant PayloadSizeInBytes : integer := PayloadSize*4;
   begin
      y(1) := x"61";
      y(2) := std_logic_vector(to_unsigned(PayloadSizeInBytes,8)); -- Payload size
      
      for i in 1 to PayloadSize loop
         case i is
            when 1  => data32_slv := std_logic_vector(resize(a.ZSIZE	   , 32));
            when 2  => data32_slv := std_logic_vector(resize(a.XSIZE	   , 32));
            when 3  => data32_slv := std_logic_vector(resize(a.YSIZE		, 32));
            when 4  => data32_slv := std_logic_vector(resize(a.IMGSIZE  , 32));
            when 5  => data32_slv := std_logic_vector(resize(a.TAGSIZE	, 32));
            when 6  => data32_slv := std_logic_vector(resize(a.SB_Min   , 32));
            when 7  => data32_slv := std_logic_vector(resize(a.SB_Max   , 32));
            when 8  => data32_slv := std_logic_vector(resize(a.SB_Mode  , 32));
            when 9  => data32_slv := std_logic_vector(resize(unsigned(a.Interleave) , 32)); 
            when 10 => data32_slv := std_logic_vector(resize(unsigned(a.Mode)       , 32));
            --when 10 => data32_slv := std_logic_vector(resize(unsigned(a.Mode) + to_unsigned(MissingImages*65536,32) , 32));
            when 11 => data32_slv := std_logic_vector(resize(a.AVGSIZE	  , 32));
            --when 12 => data32_slv := std_logic_vector(resize(a.DIAGSIZE   , 32));
            when 12 => data32_slv := std_logic_vector(resize(unsigned(a.DIAGSIZE) + to_unsigned(MissingImages*65536,32) , 32));
            when 13 => data32_slv := std_logic_vector(resize(a.BB_Temp    , 32));
            when 14 => data32_slv := std_logic_vector(resize(unsigned(a.Delta_OPD)  , 32));
            when 15 => data32_slv := std_logic_vector(resize(a.Max_Temp   , 32));
            when 16 => data32_slv := std_logic_vector(resize(a.SB_Min_Cal   , 32));
            when 17 => data32_slv := std_logic_vector(resize(a.SB_Max_Cal    , 32));
            --when 18 => data32_slv := std_logic_vector(resize(a.Lh_Exp     , 32));
            --when 19 => data32_slv := std_logic_vector(resize(a.DLbb_Exp   , 32));
         end case;
         
         y(i*4-3 + 2) := data32_slv(31 downto 24); -- MSB
         y(i*4-2 + 2) := data32_slv(23 downto 16);
         y(i*4-1 + 2) := data32_slv(15 downto 8);
         y(i*4 + 2)   := data32_slv(7 downto 0);-- LSB
      end loop;
      
      return y;
   end to_DPConfig_array8;   
   -- pragma translate_on
   
   -- pragma translate_off
   function to_DPConfig (a: DPConfig_array8) return DPConfig is
      variable y : DPConfig;
   begin
      assert FALSE report "Function not supported (probably never will)" severity FAILURE;
      return y;
   end to_DPConfig;
   
   function to_DPConfig (a: DPBConfig; Mode : std_logic_vector) return DPConfig is
      variable y : DPConfig;
   begin
      y.ZSIZE      := a.Fringe_Total;
      y.XSIZE	    := a.XSIZE;
      y.YSIZE		 := a.YSIZE;
      y.IMGSIZE    := a.IMGSIZE;
      y.TAGSIZE	 := a.TAGSIZE;
      y.SB_Min     := a.SpectralBand_Param.Min;
      y.SB_Max     := a.SpectralBand_Param.Max;
      y.SB_Mode    := unsigned(a.SpectralBand_Param.Mode);
      y.Interleave := a.Datacube_Interleave;
      
      y.Mode	    := Mode;
      y.AVGSIZE	 := a.AVGSIZE;
      y.DIAGSIZE   := x"0001";
      y.BB_Temp    := (others => '0');
      y.Delta_OPD  := (others => '0');
      y.Max_Temp   := (others => '0');
      y.SB_Min_Cal := a.SpectralBand_Param.Min;
      y.SB_Max_Cal := a.SpectralBand_Param.Max;
      --y.Lh_Exp     := (others => '0');
      --y.DLbb_Exp   := (others => '0');
      return y;
   end to_DPConfig;
   -- pragma translate_on
   
   -- pragma translate_off
   function to_DCUBE_HEADER_array (a: DPConfig; b: CLinkConfig) return DCUBE_HEADER_array is
      variable y : DCUBE_HEADER_array;
      variable Mode : std_logic_vector(7 downto 0);
   begin
      for i in 1 to 512 loop
         y(i) := x"00";
      end loop;
      
      y(1)  := x"76";
      y(2)  := x"33";
      
      -- Laser wavelength
      y(33) := x"E0";
      y(34) := x"A7";
      y(35) := x"09";
      y(36) := x"00";
      
      y(57) := x"01";
      
      Mode := ('0' & a.Mode(6 downto 0));
      if (Mode = DP_IGM or Mode = DP_HOT_BB_OUT or Mode = DP_COLD_BB_OUT) then
         y(58) := x"00"; -- Output Type : IGM
         y(59) := x"00"; -- DataFormat : UINT
      elsif (Mode = DP_RAW_SPC) then
         y(58) := x"01"; -- Output Type : RAW COMP
         y(59) := x"01"; -- DataFormat : block floating point
      elsif (Mode = DP_CAL_SPC_ONLY) then
         y(58) := x"05"; -- Output Type : SPC CAL REAL
         y(59) := x"01"; -- DataFormat : block floating point
      elsif (Mode = DP_CAL_SPC_N_IGM) then
         y(58) := x"08"; -- Output Type : IGM AND SPC CAL REAL
         y(59) := x"63"; -- DataFormat : mixed??
      elsif (Mode = DP_GAIN_OFFSET) then
         y(58) := x"07"; -- Output Type : IGM AND SPC CAL REAL
         y(59) := x"01"; -- DataFormat : block floating point
      else
         assert FALSE report "Mode not supported!!!" severity ERROR;
      end if;
      
      y(60) := x"02"; -- PixelSize
      y(61) := "000000" & a.Interleave;
      y(62) := "000000" & std_logic_vector(a.SB_Mode);
      y(63 to 66) := (std_logic_vector(a.SB_Min(7 downto 0)), std_logic_vector(a.SB_Min(15 downto 8)), x"00", x"00");
      y(67 to 70) := (std_logic_vector(a.SB_Max(7 downto 0)), std_logic_vector(a.SB_Max(15 downto 8)), x"00", x"00");
      y(71 to 72) := (std_logic_vector(b.LValSize(7 downto 0)), std_logic_vector(b.LValSize(15 downto 8)));
      y(75 to 76) := (std_logic_vector(b.HeaderSize(7 downto 0)), std_logic_vector(b.HeaderSize(15 downto 8)));
      y(77 to 78) := (std_logic_vector(a.XSIZE(7 downto 0)), "000000" & std_logic_vector(a.XSIZE(9 downto 8)));
      y(79 to 80) := (std_logic_vector(a.YSIZE(7 downto 0)), "000000" & std_logic_vector(a.YSIZE(9 downto 8)));
      y(101) := std_logic_vector(a.TAGSIZE);
      y(102) := "00" & std_logic_vector(a.AVGSIZE);
      y(136 to 139) := (std_logic_vector(a.ZSIZE(7 downto 0)), std_logic_vector(a.ZSIZE(15 downto 8)), std_logic_vector(a.ZSIZE(23 downto 16)), x"00");
      y(157) := x"04";
      y(158) := x"01";
      y(173 to 174) := (x"01", x"00"); -- BinX
      y(175 to 176) := (x"01", x"00"); -- BinY
      
      if (Mode = DP_COLD_BB_OUT) then
         y(222) := x"01";
         y(227 to 228) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
         y(229 to 230) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
      elsif (Mode = DP_HOT_BB_OUT) then
         y(222) := x"02";
         y(227 to 228) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
         y(229 to 230) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
      else
         y(222) := x"00";
      end if;
      
      return y;
   end to_DCUBE_HEADER_array;
   
   function to_DCUBE_Header_part1_array8_v4(a: DPConfig; b: CLinkConfig; SamplingPeriodNumerator: std_logic_vector) return DCUBE_Header_part1_array8_v4 is
      variable y : DCUBE_Header_part1_array8_v4; 
      variable Mode : std_logic_vector(7 downto 0);
      variable k : integer := 1;
   begin
      for i in 1 to DCUBE_Part1_V4_size loop
         y(i) := x"00";
      end loop;            
      
      y(1)  := x"76";
      y(2)  := x"34";
      k := 3;
      
      -- Laser wavelength
      y(33) := x"E0";
      y(34) := x"A7";
      y(35) := x"09";
      y(36) := x"00";      
      
      --      -- Instrument Information
      --      for i in 1 to 58  loop
      --         y(k) := x"00";
      --         k := k + 1;
      --      end loop;                      
      
      y(61) := x"01"; -- Operating Mode
      
      -- Output Type and Data Format
      Mode := ('0' & a.Mode(6 downto 0));
      if (Mode = DP_IGM or Mode = DP_HOT_BB_OUT or Mode = DP_COLD_BB_OUT) then
         y(62) := x"00"; -- Output Type : IGM
         y(63) := x"00"; -- DataFormat : UINT
      elsif (Mode = DP_RAW_SPC) then
         y(62) := x"01"; -- Output Type : RAW COMP
         y(63) := x"01"; -- DataFormat : block floating point
      elsif (Mode = DP_RAW_SPC_N_IGM) then
         y(62) := x"09"; -- Output Type : OUTPUT_TYPE_SENSOR_IGM_AND_SPC_RAW_COMP
         y(63) := x"01"; -- DataFormat : DATA_FORMAT_16B_BLOCK_FLOAT   
      elsif (Mode = DP_CAL_SPC_ONLY) then
         y(52) := x"05"; -- Output Type : SPC CAL REAL
         y(63) := x"01"; -- DataFormat : block floating point
      elsif (Mode = DP_CAL_SPC_N_IGM) then
         y(62) := x"08"; -- Output Type : IGM AND SPC CAL REAL
         y(63) := x"63"; -- DataFormat : mixed??
      elsif (Mode = DP_GAIN_OFFSET) then
         y(62) := x"07"; -- Output Type : IGM AND SPC CAL REAL
         y(63) := x"01"; -- DataFormat : block floating point
      else
         assert FALSE report "Mode not supported!!!" severity ERROR;
      end if;
      
      y(64) := x"02"; -- BytesPerPixel
      y(65) := "000000" & a.Interleave;
      y(66) := "000000" & std_logic_vector(a.SB_Mode);
      y(67 to 70) := (std_logic_vector(a.SB_Min(7 downto 0)), std_logic_vector(a.SB_Min(15 downto 8)), x"00", x"00");
      y(71 to 74) := (std_logic_vector(a.SB_Max(7 downto 0)), std_logic_vector(a.SB_Max(15 downto 8)), x"00", x"00");
      y(75 to 78) := (std_logic_vector(a.SB_Min_Cal(7 downto 0)), std_logic_vector(a.SB_Min_Cal(15 downto 8)), x"00", x"00");
      y(79 to 82) := (std_logic_vector(a.SB_Max_Cal(7 downto 0)), std_logic_vector(a.SB_Max_Cal(15 downto 8)), x"00", x"00");      
      y(83 to 86) := (std_logic_vector(a.Max_Temp(7 downto 0)), std_logic_vector(a.Max_Temp(15 downto 8)), x"00", x"00");      
      y(87 to 88) := (std_logic_vector(b.LValSize(7 downto 0)), std_logic_vector(b.LValSize(15 downto 8)));
      y(91 to 94) := (std_logic_vector(b.HeaderSize(7 downto 0)), std_logic_vector(b.HeaderSize(15 downto 8)), x"00", x"00");
      y(95 to 96) := (std_logic_vector(a.XSIZE(7 downto 0)), "000000" & std_logic_vector(a.XSIZE(9 downto 8)));
      y(97 to 98) := (std_logic_vector(a.YSIZE(7 downto 0)), "000000" & std_logic_vector(a.YSIZE(9 downto 8)));
      y(119) := std_logic_vector(a.TAGSIZE);
      y(120) := "00" & std_logic_vector(a.AVGSIZE);
      y(165 to 168) := (std_logic_vector(a.ZSIZE(7 downto 0)), std_logic_vector(a.ZSIZE(15 downto 8)), std_logic_vector(a.ZSIZE(23 downto 16)), x"00");   
      y(186) := SamplingPeriodNumerator; -- SamplingPeriodNumerator
      y(187) := x"01"; -- SamplingPeriodDenominator
      y(202 to 203) := (x"01", x"00"); -- BinX
      y(204 to 205) := (x"01", x"00"); -- BinY
      
      if (Mode = DP_COLD_BB_OUT) then
         y(280) := x"01"; -- InputBB
         y(285 to 286) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
         y(287 to 288) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
      elsif (Mode = DP_HOT_BB_OUT) then
         y(280) := x"02";
         y(285 to 286) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
         y(287 to 288) :=  (std_logic_vector(a.BB_Temp(7 downto 0)), std_logic_vector(a.BB_Temp(15 downto 8)));
      else
         y(280) := x"00";
      end if;
      
      return y;
   end to_DCUBE_Header_part1_array8_v4;
   
   -- pragma translate_on
   
   
   function to_output_debug(a: std_logic_vector(15 downto 0)) return t_output_debug is
      variable y: t_output_debug;
   begin
      y.FPGA_ID := a(15);
      y.Z := a(14 downto 10);
      y.Y := a(9 downto 5);
      y.X := a(4 downto 0);
      return y;
   end to_output_debug;
   
   
   function to_output_debug32(a: std_logic_vector(31 downto 0)) return t_output_debug32 is
      variable y: t_output_debug32;
   begin
      y.H :=to_output_debug(a(31 downto 16));
      y.L :=to_output_debug(a(15 downto 0));
      return y;
   end to_output_debug32;
   
   
   function to_ddr_data21_debug(a: std_logic_vector(127 downto 0)) return t_ddr_data21_debug is
      variable y: t_ddr_data21_debug;
   begin
      y.P0 := a(20 downto 0);
      y.P1 := a(41 downto 21);
      y.P2 := a(62 downto 42);
      y.P3 := a(83 downto 63);
      y.P4 := a(104 downto 84);
      y.P5 := a(125 downto 105);
      return y;
   end to_ddr_data21_debug;
   
   function to_std_logic_vector (a: VP30StatusInfo) return std_logic_vector is
      variable y: std_logic_vector(47 downto 0);
   begin
      y(47 downto 40) := a.ExtTemp;
      y(39 downto 32) := a.IntTemp;
      y(31 downto 0)  := a.Stat;
      return y;
   end to_std_logic_vector;
   
   function to_VP30StatusInfo (a: std_logic_vector) return VP30StatusInfo is
      variable y: VP30StatusInfo;
   begin
      y.ExtTemp := a(47 downto 40);
      y.IntTemp := a(39 downto 32);
      y.Stat    := a(31 downto 0);
      return y;
   end to_VP30StatusInfo;
   
   function to_std_logic_vector (a: VP7StatusInfo) return std_logic_vector is
      variable y: std_logic_vector(47 downto 0);
   begin
      y(47 downto 40) := a.ExtTemp;
      y(39 downto 32) := a.IntTemp;
      y(31 downto 0)  := a.Stat;
      return y;
   end to_std_logic_vector;
   
   function to_VP7StatusInfo (a: std_logic_vector) return VP7StatusInfo is
      variable y: VP7StatusInfo;
      
   begin
      y.ExtTemp := a(47 downto 40);
      y.IntTemp := a(39 downto 32);
      y.Stat    := a(31 downto 0);
      return y;
   end to_VP7StatusInfo;
   
   function status_latch (new_status,old_status: VP30StatusInfo) return VP30StatusInfo is
      variable y : VP30StatusInfo;
   begin
      y.ExtTemp            := Uto0(new_status.ExtTemp);
      y.IntTemp            := Uto0(new_status.IntTemp);
      
      -- Latch all bits
      y.Stat               := Uto0(old_status.Stat) or Uto0(new_status.Stat);
      
      -- Renew only certain bits (which are not error bits)
      y.Stat(2)            := Uto0(new_status.Stat)(2);
      y.Stat(9 downto 8)   := Uto0(new_status.Stat)(9 downto 8);
      y.Stat(11)           := Uto0(new_status.Stat)(11);
      
      return y;
   end status_latch;
   
   function status_latch (new_status,old_status: VP7StatusInfo) return VP7StatusInfo is
      variable y : VP7StatusInfo;
   begin
      y.ExtTemp            := Uto0(new_status.ExtTemp);
      y.IntTemp            := Uto0(new_status.IntTemp);
      y.Stat               := Uto0(new_status.Stat) or Uto0(old_status.Stat);
      return y;
   end status_latch;            
   
   function to_ROIC_CLink_Header_array16(h: ROIC_DCube_Header; f: ROIC_DCube_Footer) return ROIC_CLink_Header_array16 is
      variable y: ROIC_CLink_Header_array16;
   begin
      y(1)  := x"00" & h.Direction & std_logic_vector(h.Acq_Number(22 downto 16));
      y(2)  := std_logic_vector(h.Acq_Number(15 downto 0));
      y(3)  := x"00" & std_logic_vector(f.Write_No(23 downto 16));
      y(4)  := std_logic_vector(f.Write_No(15 downto 0));
      y(5)  := x"00" & std_logic_vector(f.Trig_No(23 downto 16));
      y(6)  := std_logic_vector(f.Trig_No(15 downto 0));
      y(7)  := std_logic_vector(h.Code_Rev);
      --y(8)  := x"0000"; -- SpareA
      y(8)  := std_logic_vector(f.Status(31 downto 16));
      y(9)  := std_logic_vector(f.Status(15 downto 0));
      y(10)  := (15 downto RXLEN => '0') & std_logic_vector(h.Xmin);
      y(11) := (15 downto RYLEN => '0') & std_logic_vector(h.Ymin);
      y(12) := x"00" & std_logic_vector(f.ZPDPosition(23 downto 16));
      y(13) := std_logic_vector(f.ZPDPosition(15 downto 0));
      y(14) := std_logic_vector(f.ZPDPeakVal);
      y(15) := std_logic_vector(h.StartTimeStamp(31 downto 16));
      y(16) := std_logic_vector(h.StartTimeStamp(15 downto 0));
      y(17) := std_logic_vector(f.EndTimeStamp(31 downto 16));
      y(18) := std_logic_vector(f.EndTimeStamp(15 downto 0));      
      return y;
   end to_ROIC_CLink_Header_array16; 
   
   function to_ROIC_CLink_Header_array16_v4(h: ROIC_DCube_Header_v2_6;f: ROIC_DCube_Footer_v2_6; DP_Present :std_logic) return ROIC_CLink_Header_array16_v4 is
      variable y: ROIC_CLink_Header_array16_v4;
   begin 
      if DP_Present= '1' then         
         -- footer status
         y(1)  := std_logic_vector(f.Status(31 downto 16));       
         y(2)  := std_logic_vector(f.Status(15 downto 0));          
      else  -- then Clink connected to Roic
         -- header status
         y(1)  := std_logic_vector(h.Status(31 downto 16));       
         y(2)  := std_logic_vector(h.Status(15 downto 0));   
      end if;
      -- ROIC_header part
      y(3)  := x"00" & h.Direction & std_logic_vector(h.Acq_Number(22 downto 16)); 
      y(4)  := std_logic_vector(h.Acq_Number(15 downto 0)); 
      y(5)  := x"0000";  -- code revision MSB 16 bits
      y(6)  := std_logic_vector(h.Code_Rev);
      y(7)  := (15 downto RXLEN => '0') & std_logic_vector(h.Xmin);
      y(8)  := (15 downto RYLEN => '0') & std_logic_vector(h.Ymin); 
      y(9)  := std_logic_vector(h.StartTimeStamp(31 downto 16));
      y(10) := std_logic_vector(h.StartTimeStamp(15 downto 0));
      y(11) := std_logic_vector(resize(h.FPGATemp,16));
      y(12) := std_logic_vector(resize(h.PCBTemp,16));
      y(13) := (15 downto 2 => '0') & h.FilterPosition;
      y(14) := (15 downto 1 => '0') & std_logic(h.ArmedStatus);        
      y(15) := std_logic_vector(h.RealIntTime);    
      y(16) := std_logic_vector(h.Spare); 
      if DP_Present= '1' then
         -- ROIC_Footer part
         y(17) := x"0000";
         y(18) := std_logic_vector(f.Write_No(15 downto 0));
         y(19) := x"0000";
         y(20) := std_logic_vector(f.Trig_No(15 downto 0));
         y(21) := x"0000";
         y(22) := std_logic_vector(f.ZPDPosition(15 downto 0));
         y(23) := x"0000";
         y(24) := std_logic_vector(f.ZPDPeakVal(15 downto 0));
         y(25) := std_logic_vector(f.EndTimeStamp(31 downto 16));
         y(26) := std_logic_vector(f.EndTimeStamp(15 downto 0)); 
         y(27) := std_logic_vector(f.NbPixelsAboveHighLimit(31 downto 16));
         y(28) := std_logic_vector(f.NbPixelsAboveHighLimit(15 downto 0)); 
         y(29) := std_logic_vector(f.NbPixelsAboveLowLimit(31 downto 16));
         y(30) := std_logic_vector(f.NbPixelsAboveLowLimit(15 downto 0)); 
         y(31) := f.Nav_Data_Tag(31 downto 16);
         y(32) := f.Nav_Data_Tag(15 downto 0); 
      else
         for i in 17 to 32 loop
            y(i) := (others => '0');
         end loop;
      end if;
      return y;
   end to_ROIC_CLink_Header_array16_v4;  
   
   function to_NAV_CLINK_Header_array16_v4(h: NAV_DCube_Header_v2_6) return NAV_CLINK_Header_array16_v4 is
      variable y: NAV_CLINK_Header_array16_v4;
   begin 
      for i in  1 to NAV_DATA_REAL_V4_SIZE/4 loop
         y(2*i-1)  := h(i)(31 downto 16);
         y(2*i):= h(i)(15 downto 0);
      end loop;      
      return y;
   end to_NAV_CLINK_Header_array16_v4;
   
   function to_ROIC_CLink_Header_array16(h: ROIC_DCube_Header) return ROIC_CLink_Header_array16 is
      variable y: ROIC_CLink_Header_array16;
   begin
      y(1)  := x"00" & h.Direction & std_logic_vector(h.Acq_Number(22 downto 16));
      y(2)  := std_logic_vector(h.Acq_Number(15 downto 0));
      y(3)  := x"0000";
      y(4)  := x"0000";
      y(5)  := x"0000";
      y(6)  := x"0000";
      y(7)  := std_logic_vector(h.Code_Rev);
      --y(8)  := x"0000"; -- SpareA
      y(8)  := std_logic_vector(h.Status(31 downto 16));
      y(9)  := std_logic_vector(h.Status(15 downto 0));
      y(10)  := (15 downto RXLEN => '0') & std_logic_vector(h.Xmin);
      y(11) := (15 downto RYLEN => '0') & std_logic_vector(h.Ymin);
      y(12) := x"0000";
      y(13) := x"0000";
      y(14) := x"0000";
      y(15) := std_logic_vector(h.StartTimeStamp(31 downto 16));
      y(16) := std_logic_vector(h.StartTimeStamp(15 downto 0));
      y(17) := x"0000";
      y(18) := x"0000";
      return y;
   end to_ROIC_CLink_Header_array16;  
   
   --function to_ROIC_CLink_Header_array16_v4(h: ROIC_DCube_Header_v2_6) return ROIC_CLink_Header_array16_v4 is
   --   variable y: ROIC_CLink_Header_array16_v4;
   --begin
   --   y(1)  := std_logic_vector(h.Status(31 downto 16));
   --   y(2)  := std_logic_vector(h.Status(15 downto 0));
   --   y(3)  := x"00" & h.Direction & std_logic_vector(h.Acq_Number(22 downto 16)); 
   --   y(4)  := std_logic_vector(h.Acq_Number(15 downto 0)); 
   --   y(5)  := x"0000";  -- code revision MSB 16 bits
   --   y(6)  := std_logic_vector(h.Code_Rev);
   --   y(7)  := (15 downto RXLEN => '0') & std_logic_vector(h.Xmin);
   --   y(8)  := (15 downto RYLEN => '0') & std_logic_vector(h.Ymin); 
   --   y(9)  := std_logic_vector(h.StartTimeStamp(31 downto 16));
   --   y(10) := std_logic_vector(h.StartTimeStamp(15 downto 0));
   --   
   --   y(11) := std_logic_vector(resize(h.FPGATemp,16));
   --   y(12) := std_logic_vector(resize(h.PCBTemp,16));
   --   y(13) := (15 downto 1 => '0') & std_logic(h.FilterPosition);
   --   y(14) := (15 downto 1 => '0') & std_logic(h.ArmedStatus);        
   --   y(15) := std_logic_vector(h.RealIntTime);    
   --   y(16) := std_logic_vector(h.Spare); 
   --   -- ROIC_Footer part ( non existant)
   --   y(17) := x"0000";
   --   y(18) := x"0000";
   --   y(19) := x"0000";
   --   y(20) := x"0000";     
   --   y(21) := x"0000";
   --   y(22) := x"0000";
   --   y(23) := x"0000";      
   --   y(24) := x"0000";
   --   y(25) := x"0000";
   --   y(26) := x"0000";      
   --   y(27) := x"0000";
   --   y(28) := x"0000";
   --   y(29) := x"0000";
   --   y(30) := x"0000";     
   --   y(31) := x"0000";
   --   y(32) := x"0000";
   --   
   --   return y;
   --end to_ROIC_CLink_Header_array16_v4;
   
   
   function to_DCUBE_FOOTER_V3_array (a, b : DPB_DCube_Header; c : VP7StatusInfo) return DCUBE_FOOTER_V3_array is
      variable y: DCUBE_FOOTER_V3_array;
      --variable ROICInfo: ROIC_Img_Footer;
      variable ROICInfo_ary: ROIC_CLink_Header_array16;
   begin
      -- ROIC Section (1 to 18)
      --      ROICInfo := to_ROIC_Img_Footer(a.ROICHeader, a.ROICFooter);
      --      ROICInfo_ary := to_ROIC_Img_Footer_array16(ROICInfo);
      ROICInfo_ary := to_ROIC_CLink_Header_array16(a.ROICHeader, a.ROICFooter);
      for i in ROICInfo_ary'range loop
         y(i) := ROICInfo_ary(i);
      end loop;
      
      -- DPB Section (17 to 44)
      --y(17) := x"0000";                                                   -- SpareB
      --y(18) := x"0000";                                                   -- SpareB
      y(19) := a.VP30Status.Stat(31 downto 16);
      y(20) := a.VP30Status.Stat(15 downto 0);
      y(21) := a.VP30Status.IntTemp & a.VP30Status.ExtTemp;           -- DCA_FPGA1_Temp & FPGA1_ExtTemp
      y(22) := X"0000";                                                  -- Spare C
      y(23) := x"0000";                                                  -- Spare C
      y(24) := b.VP30Status.Stat(31 downto 16);
      y(25) := b.VP30Status.Stat(15 downto 0);
      y(26) := b.VP30Status.IntTemp & b.VP30Status.ExtTemp;           -- DCA_FPGA2_Temp & FPGA2_ExtTemp
      y(27) := X"0000";                                                  -- Spare D
      y(28) := X"0000";                                                  -- Spare D
      y(29) := c.Stat(31 downto 16);
      y(30) := c.Stat(15 downto 0);
      y(31) := c.IntTemp & c.ExtTemp;                                 -- DCA_FPGA3_Temp & FPGA3_ExtTemp
      y(32) := "000" & std_logic_vector(a.DUI(28 downto 16));            -- DCA_DUI hi
      y(33) := std_logic_vector(a.DUI(15 downto 0));                     -- DCA_DUI lo
      y(34) := X"0000";                                      -- DCA_DPBFirmwareVersion
      y(35) := X"0000";                                                  -- Spare E
      y(36) := X"0000";                                                  -- Spare E
      y(37) := X"0000";                                                  -- Spare E
      y(38) := X"0000";                                                  -- Spare E
      y(39) := X"0000";                                                  -- Spare E
      y(40) := X"0000";                                                  -- Spare E
      y(41) := X"0000";                                                  -- Spare E
      y(42) := X"0000";                                                  -- Spare E
      y(43) := X"0000";                                                  -- Spare E
      y(44) := X"0000";                                                  -- Spare E
      
      return y;
   end to_DCUBE_FOOTER_V3_array;
   
   function to_DCUBE_Header_Part2_array_V4 (a, b : DPB_DCube_Header_v2_6; c : VP7StatusInfo; DP_Present:Std_logic) return DCUBE_Header_Part2_array_V4 is
      variable y : DCUBE_Header_Part2_array_V4;
      variable DP1 : DPB_DCube_Header_array32_v2_6;
      variable DP2 : DPB_DCube_Header_array32_v2_6;
      variable ROICInfo_ary: ROIC_CLink_Header_array16_v4;
      variable NAVInfo_ary: NAV_CLink_Header_array16_v4;
      variable k : integer := 1;
   begin
      -- Roic part------------------------------------------------
      ROICInfo_ary := to_ROIC_CLink_Header_array16_v4(a.ROICHeader, a.ROICFooter, DP_Present);
      for i in ROICInfo_ary'range loop
         y(k) := ROICInfo_ary(i); 
         k := k + 1;
      end loop; 
      
      -- SpareA_V4
      for i in 1 to SPAREA_LEN_V4/2  loop
         y(k) := x"AAAA";
         k := k + 1;
      end loop; 
      
      -- Geopositionning part--------------------------------------
      --      for i in 1 to GEOPOS_LEN_V4/2 loop
      --         y(k) := (others =>'0');
      --         k := k + 1;
      --      end loop; 
      NAVInfo_ary := to_NAV_CLINK_Header_array16_v4(a.NAVHeader);
      for i in NAVInfo_ary'range loop
         y(k) := NAVInfo_ary(i); 
         k := k + 1;
      end loop; 
      
      -- SpareB_V4
      if SPAREB_LEN_V4 > 2 then  
         for i in 1 to SPAREB_LEN_V4/2  loop
            y(k) := x"BBBB";
            k := k + 1;
         end loop; 
      end if;
      -- DPB part---------------------------------------------------         
      
      -- SpareC
      for i in 1 to SPAREC_LEN_V4/2  loop
         y(k) := x"CCCC";
         k := k + 1;
      end loop; 
      
      if DP_Present = '1' then
         DP1 := to_DPB_DCube_Header_array32_v2_6(a);      
         for i in 2 to DPB_DCube_Header_v2_6_32_LEN  loop
            y(k) := DP1(i)(31 downto 16);
            k := k + 1;
            y(k) := DP1(i)(15 downto 0); 
            k := k + 1;
         end loop;     
      else
         for i in 2 to DPB_DCube_Header_v2_6_32_LEN  loop
            y(k) := (others => '0');
            k := k + 1;
            y(k) := (others => '0');
            k := k + 1;
         end loop;        
      end if;
      
      -- SpareD
      for i in 1 to SPARED_LEN_V4/2  loop
         y(k) := x"DDDD";   
         k := k + 1;
      end loop;
      
      if DP_Present = '1' then
         DP2 := to_DPB_DCube_Header_array32_v2_6(b);  
         for i in 2 to DPB_DCube_Header_v2_6_32_LEN  loop
            y(k) := DP2(i)(31 downto 16);
            k := k + 1;
            y(k) := DP2(i)(15 downto 0); 
            k := k + 1;
         end loop;   
      else
         for i in 2 to DPB_DCube_Header_v2_6_32_LEN  loop
            y(k) := (others => '0');
            k := k + 1;
            y(k) := (others => '0');
            k := k + 1;
         end loop;        
      end if;           
      
      -- SpareE
      for i in 1 to SPAREE_LEN_V4/2  loop
         y(k) := x"EEEE";  
         k := k + 1;
      end loop;
      
      
      --CLINK info---------------------------------------------------------------
      y(k) := c.Stat(31 downto 16);   
      k := k + 1;
      y(k) := c.Stat(15 downto 0);  
      k := k + 1;
      y(k) := c.IntTemp & c.ExtTemp;
      k := k + 1;
      y(k) := std_logic_vector(resize(unsigned(CLINK_VERSION),y(k)'LENGTH));
      k := k + 1;  
      
      -- SpareF
      for i in 1 to SPAREF_LEN_V4/2  loop
         y(k) := x"FFFF";
         k := k + 1;
      end loop;
      
      assert (k = DCUBE_Header_Part2_array_V4'LENGTH+1) report "DCUBE_Header_Part2_array_V4 was not assigned properly!" severity FAILURE;
      
      return y;
   end to_DCUBE_Header_Part2_array_V4;   
   
   
   
   function to_DCUBE_FOOTER_V3_array (a: ROIC_DCube_Header; c : VP7StatusInfo) return DCUBE_FOOTER_V3_array is
      variable y: DCUBE_FOOTER_V3_array;
      --variable ROICInfo: ROIC_Img_Footer;
      variable ROICInfo_ary: ROIC_CLink_Header_array16;
   begin
      -- ROIC Section (1 to 18)
      --      ROICInfo := to_ROIC_Img_Footer(a.ROICHeader, a.ROICFooter);
      --      ROICInfo_ary := to_ROIC_Img_Footer_array16(ROICInfo);
      ROICInfo_ary := to_ROIC_CLink_Header_array16(a);
      for i in ROICInfo_ary'range loop
         y(i) := ROICInfo_ary(i);
      end loop;
      
      -- DPB Section (17 to 44)
      --y(17) := x"0000";                -- SpareB
      --y(18) := x"0000";                -- SpareB
      y(19) := x"0000";
      y(20) := x"0000";
      y(21) := x"0000";                -- DCA_FPGA1_Temp & FPGA1_ExtTemp
      y(22) := X"0000";                -- Spare C
      y(23) := x"0000";                -- Spare C
      y(24) := x"0000";
      y(25) := x"0000";
      y(26) := x"0000";                -- DCA_FPGA2_Temp & FPGA2_ExtTemp
      y(27) := X"0000";                -- Spare D
      y(28) := X"0000";                -- Spare D
      y(29) := c.Stat(31 downto 16);
      y(30) := c.Stat(15 downto 0);
      y(31) := c.IntTemp & c.ExtTemp;  -- DCA_FPGA3_Temp & FPGA3_ExtTemp
      y(32) := x"0000";                -- DCA_DUI hi
      y(33) := x"0000";                -- DCA_DUI lo
      y(34) := x"0000";                -- DCA_DPBFirmwareVersion
      y(35) := X"0000";                -- Spare E
      y(36) := X"0000";                -- Spare E
      y(37) := X"0000";                -- Spare E
      y(38) := X"0000";                -- Spare E
      y(39) := X"0000";                -- Spare E
      y(40) := X"0000";                -- Spare E
      y(41) := X"0000";                -- Spare E
      y(42) := X"0000";                -- Spare E
      y(43) := X"0000";                -- Spare E
      y(44) := X"0000";                -- Spare E
      
      return y;
   end to_DCUBE_FOOTER_V3_array;
   
   --function to_DCUBE_Part2_V4_array (a: ROIC_DCube_Header_v2_6; c : VP7StatusInfo) return DCUBE_Part2_V4_array is
   --      variable y: DCUBE_Part2_V4_array;
   --      --variable ROICInfo: ROIC_Img_Footer;
   --      variable ROICInfo_ary: ROIC_CLink_Header_array16;
   --   begin
   --      -- ROIC Section (1 to 18)
   --      --      ROICInfo := to_ROIC_Img_Footer(a.ROICHeader, a.ROICFooter);
   --      --      ROICInfo_ary := to_ROIC_Img_Footer_array16(ROICInfo);
   --      ROICInfo_ary := to_ROIC_CLink_Header_array16(a);
   --      for i in ROICInfo_ary'range loop
   --         y(i) := ROICInfo_ary(i);
   --      end loop;
   --      
   --      -- DPB Section (17 to 44)
   --      --y(17) := x"0000";                -- SpareB
   --      --y(18) := x"0000";                -- SpareB
   --      y(19) := x"0000";
   --      y(20) := x"0000";
   --      y(21) := x"0000";                -- DCA_FPGA1_Temp & FPGA1_ExtTemp
   --      y(22) := X"0000";                -- Spare C
   --      y(23) := x"0000";                -- Spare C
   --      y(24) := x"0000";
   --      y(25) := x"0000";
   --      y(26) := x"0000";                -- DCA_FPGA2_Temp & FPGA2_ExtTemp
   --      y(27) := X"0000";                -- Spare D
   --      y(28) := X"0000";                -- Spare D
   --      y(29) := c.Stat(31 downto 16);
   --      y(30) := c.Stat(15 downto 0);
   --      y(31) := c.IntTemp & c.ExtTemp;  -- DCA_FPGA3_Temp & FPGA3_ExtTemp
   --      y(32) := x"0000";                -- DCA_DUI hi
   --      y(33) := x"0000";                -- DCA_DUI lo
   --      y(34) := x"0000";                -- DCA_DPBFirmwareVersion
   --      y(35) := X"0000";                -- Spare E
   --      y(36) := X"0000";                -- Spare E
   --      y(37) := X"0000";                -- Spare E
   --      y(38) := X"0000";                -- Spare E
   --      y(39) := X"0000";                -- Spare E
   --      y(40) := X"0000";                -- Spare E
   --      y(41) := X"0000";                -- Spare E
   --      y(42) := X"0000";                -- Spare E
   --      y(43) := X"0000";                -- Spare E
   --      y(44) := X"0000";                -- Spare E
   --      
   --      return y;
   --   end to_DCUBE_Part2_V4_array;
   
   function to_DCUBE_FOOTER_V3 (b: DCUBE_FOOTER_V3_array) return DCUBE_FOOTER_V3 is
      variable a : DCUBE_FOOTER_V3_array8;
      variable y: DCUBE_FOOTER_V3;
      variable Stat1 : std_logic_vector(47 downto 0);
      variable Stat2 : std_logic_vector(47 downto 0);
      variable Stat3 : std_logic_vector(47 downto 0);
      
   begin
      for i in DCUBE_FOOTER_V3_array'range loop
         a(i*2-1) := b(i)(15 downto 8);
         a(i*2) := b(i)(7 downto 0);
      end loop;
      --y.Unused1                  := a(1);
      y.DCA_SweepDirection       := a(2)(7);
      y.DCA_DataCubeID           := unsigned(a(2)(6 downto 0)) & unsigned(a(3)) & unsigned(a(4));
      y.DCA_IntFramesCnt         := unsigned(a(5)) & unsigned(a(6)) & unsigned(a(7)) & unsigned(a(8));
      y.DCA_SampTrigsCnt         := unsigned(a(9)) & unsigned(a(10)) & unsigned(a(11)) & unsigned(a(12));
      y.DCA_ROICFirmwareVersion  := a(13) & a(14);
      --y.SpareA                   := a(15) & a(16);
      y.DCA_ROICStatus           := a(16) & a(18);
      y.DCA_FOVStartX            := unsigned(a(19)) & unsigned(a(20));
      y.DCA_FOVStartY            := unsigned(a(21)) & unsigned(a(22));
      y.DCA_ZPDPosition          := unsigned(a(23)) & unsigned(a(24)) & unsigned(a(25)) & unsigned(a(26));
      y.DCA_MaxFPACount          := unsigned(a(27)) & unsigned(a(28));
      y.DCA_TimeStamp            := unsigned(a(29)) & unsigned(a(30)) & unsigned(a(31)) & unsigned(a(32));
      --y.SpareB                   := a(33) & a(34) & a(35) & a(36);
      --y.Unused2                  := a(37);
      Stat1                      := a(42) & a(41) & b(19) & b(20);
      y.DCA_FPGA1_Status         := to_VP30StatusInfo(Stat1);
      --y.SpareC                   := a(43) & a(44) & a(45) & a(46);
      --y.Unused3                  := a(47);
      Stat2                      := a(52) & a(51) & b(24) & b(25);
      y.DCA_FPGA2_Status         := to_VP30StatusInfo(Stat2);
      --y.SpareD                   := a(53) & a(54) & a(55) & a(56);
      --y.Unused4                  := a(57);
      Stat3                      := a(62) & a(61) & b(29) & b(30);
      y.DCA_FPGA3_Status         := to_VP7StatusInfo(Stat3);
      y.DCA_DUI                  := unsigned(a(63)) & unsigned(a(64)) & unsigned(a(65)) & unsigned(a(66));
      y.DCA_DPBFirmwareVersion   := a(67) & a(68);
      --y.SpareE                  :=
      return y;
   end to_DCUBE_FOOTER_V3;
   
   -- function to_DCUBE_Header_part2_V4 (b: DCUBE_Header_part2_array_v4) return DCUBE_Header_part2_V4 is
   --      variable a : DCUBE_Header_part2_array8_v4;
   --      variable y: DCUBE_Header_part2_V4;
   --      variable Stat1 : std_logic_vector(47 downto 0);
   --      variable Stat2 : std_logic_vector(47 downto 0);
   --      variable Stat3 : std_logic_vector(47 downto 0);
   --      
   --   begin
   --      for i in DCUBE_Header_part2_array_v4'range loop
   --         a(i*2-1) := b(i)(15 downto 8);
   --         a(i*2) := b(i)(7 downto 0);
   --      end loop;                                   
   --      
   --      
   --      y.DCA_ROICStatus           := a(1) & a(2) & a(3) & a(4);
   --      y.DCA_SweepDirection       := a(6)(7);
   --      y.DCA_DataCubeID           := unsigned(a(6)(6 downto 0)) & unsigned(a(7)) & unsigned(a(8)); 
   --      y.DCA_ROICFirmwareVersion  := a(9) & a(10) & a(11) & a(12);
   --      y.DCA_FOVStartX            := unsigned(a(13)) & unsigned(a(14));
   --      y.DCA_FOVStartY            := unsigned(a(15)) & unsigned(a(16));
   --      y.DCA_Start_TimeStamp      := unsigned(a(17)) & unsigned(a(18)) & unsigned(a(19)) & unsigned(a(20));      
   --      y.DCA_ROIC_FPGATemp        := a(21) & a(22) & a(23) & a(12); 
   --      y.DCA_ROIC_FPGATemp        := a(9) & a(10) & a(11) & a(12);      
   --      y.DCA_IntFramesCnt         := unsigned(a(5)) & unsigned(a(6)) & unsigned(a(7)) & unsigned(a(8));
   --      y.DCA_SampTrigsCnt         := unsigned(a(9)) & unsigned(a(10)) & unsigned(a(11)) & unsigned(a(12));
   --      
   --      --y.SpareA                   := a(15) & a(16);
   --      
   --      
   --      y.DCA_ZPDPosition          := unsigned(a(23)) & unsigned(a(24)) & unsigned(a(25)) & unsigned(a(26));
   --      y.DCA_MaxFPACount          := unsigned(a(27)) & unsigned(a(28));
   --      
   --      --y.SpareB                   := a(33) & a(34) & a(35) & a(36);
   --      --y.Unused2                  := a(37);
   --      Stat1                      := a(42) & a(41) & b(19) & b(20);
   --      y.DCA_FPGA1_Status         := to_VP30StatusInfo(Stat1);
   --      --y.SpareC                   := a(43) & a(44) & a(45) & a(46);
   --      --y.Unused3                  := a(47);
   --      Stat2                      := a(52) & a(51) & b(24) & b(25);
   --      y.DCA_FPGA2_Status         := to_VP30StatusInfo(Stat2);
   --      --y.SpareD                   := a(53) & a(54) & a(55) & a(56);
   --      --y.Unused4                  := a(57);
   --      Stat3                      := a(62) & a(61) & b(29) & b(30);
   --      y.DCA_FPGA3_Status         := to_VP7StatusInfo(Stat3);
   --      y.DCA_DUI                  := unsigned(a(63)) & unsigned(a(64)) & unsigned(a(65)) & unsigned(a(66));
   --      y.DCA_DPBFirmwareVersion   := a(67) & a(68);
   --      --y.SpareE                  :=    
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      
   --      return y;
   --   end to_DCUBE_Header_part2_V4;
   
   function to_DPB_DCube_Header(a: unsigned(DUILEN-1 downto 0); b: VP30StatusInfo; c: ROIC_DCube_Header; d: ROIC_DCube_Footer) return DPB_DCube_Header is
      variable y : DPB_DCube_Header;
   begin
      y.DUI := a;
      y.VP30Status := b;
      y.ROICHeader := c;
      y.ROICFooter := d;
      return y;
   end to_DPB_DCube_Header;
   
   function to_DPB_DCube_Header(a: DPB_DCube_Header_array16) return DPB_DCube_Header is
      variable y : DPB_DCube_Header;
      variable stat_vec : std_logic_vector(47 downto 0);
      variable head_array : ROIC_DCube_Header_array16;
      variable foot_array : ROIC_DCube_Footer_array16;
   begin
      y.DUI := resize(unsigned(a(1)) & unsigned(a(2)), DUILEN);
      --a(3) unused
      stat_vec := a(4) & a(5) & a(6);
      y.VP30Status := to_VP30StatusInfo(stat_vec);
      
      for i in ROIC_DCube_Header_array16'range loop
         head_array(i) := a(i+6);
      end loop;
      y.ROICHeader := to_ROIC_DCube_Header(head_array);
      
      for i in ROIC_DCube_Footer_array16'range loop
         foot_array(i) := a(i+6+ROIC_DCube_Header_array16'LENGTH);
      end loop;
      y.ROICFooter := to_ROIC_DCube_Footer(foot_array);
      
      return y;
   end to_DPB_DCube_Header;
   
   function to_DPB_DCube_Header(a: DPB_DCube_Header_array32) return DPB_DCube_Header is
      variable y : DPB_DCube_Header;
      variable y1: ROIC_DCube_Header_array32;
      variable y2: ROIC_DCube_Footer_array32;
   begin
      -- SKIP Header section
      -- DPB Section
      y.DUI := unsigned(a(2)(DUILEN-1 downto 0));
      y.VP30Status.ExtTemp := a(3)(15 downto 8);
      y.VP30Status.IntTemp := a(3)(7 downto 0);
      y.VP30Status.Stat := a(4);
      -- ROIC Header Section (skip header word)
      for i in 2 to y1'length loop
         y1(i) := a(i+3);
      end loop;
      y.ROICHeader := to_ROIC_DCube_Header(y1);
      -- ROIC Footer Section (skip header word)
      for i in 2 to y2'length loop
         y2(i) := a(i+2+y1'length);
      end loop;
      y.ROICFooter := to_ROIC_DCube_Footer(y2);
      return y;
   end to_DPB_DCube_Header; 
   
   function to_DPB_DCube_Header_v2_6(a: DPB_DCube_Header_array32_v2_6) return DPB_DCube_Header_v2_6 is
      variable y : DPB_DCube_Header_v2_6;
      variable y1: ROIC_DCube_Header_array32_v2_6;
      variable y2: ROIC_DCube_Footer_array32_v2_6;
   begin
      -- DPB Section
      -- a(1), the header, is ignored.   
      y.DPBStatus         := a(2) & a(3);
      y.FirmwareVersion   := a(4)(31 downto 16);
      y.FPGATemp          := a(4)(15 downto 8);
      y.PCBTemp           := a(4)(7 downto 0);
      y.PixelsReceivedCnt := unsigned(a(5)(DUILEN-1 downto 0)); -- 4 bytes allocated for that field                     
      
      -- ROIC Header Section
      for i in 1 to y1'length loop
         y1(i) := a(i+DPB_DCube_Header_v2_6_32_LEN);
      end loop;
      y.ROICHeader := to_ROIC_DCube_Header_v2_6(y1);
      
      -- ROIC Footer Section
      for i in 1 to y2'length loop
         y2(i) := a(i+y1'length+DPB_DCube_Header_v2_6_32_LEN);
      end loop;            
      y.ROICFooter := to_ROIC_DCube_Footer_v2_6(y2); 

      -- NAV Footer Section
      for i in 1 to y.NAVHeader'length loop
         y.NAVHeader(i) := a(i+DPB_DCube_Header_v2_6_32_LEN+y1'length+y2'length);
      end loop;

      return y;
   end to_DPB_DCube_Header_v2_6;
   
   function to_DPB_DCube_Header_array32_v2_6(a: DPB_DCube_Header_v2_6) return DPB_DCube_Header_array32_v2_6 is
      variable y: DPB_DCube_Header_array32_v2_6;
      variable y1: ROIC_DCube_Header_array32_v2_6;
      variable y2: ROIC_DCube_Footer_array32_v2_6;
      variable k : integer := 1;
   begin
      -- DPB Section
      y(1) := PROC_HEADER_FRAME & std_logic_vector(to_unsigned(DPB_DCube_Header_array32_v2_6'length-1, 24)); -- Command Header + payload size
      y(2) := std_logic_vector(resize(unsigned(a.DPBStatus(DPBSTATLEN-1 downto 32)),32));
      y(3) := a.DPBStatus(31 downto 0);
      y(4) := a.FirmwareVersion & a.FPGATemp & a.PCBTemp;
      y(5) := std_logic_vector(resize(unsigned(a.PixelsReceivedCnt(DUILEN-1 downto 0)),32)); 
      k := 6;
      
      -- ROIC Header Section
      y1 := to_ROIC_DCube_Header_array32_v2_6(a.ROICHeader);     
      for i in y1'range loop
         y(k) := y1(i);  
         k := k + 1;
      end loop;
      
      -- ROIC Footer Section
      y2 := to_ROIC_DCube_Footer_array32_v2_6(a.ROICFooter);
      for i in y2'range loop
         y(k) := y2(i);  
         k := k + 1;
      end loop;
      
      -- NAV Footer Section
      for i in 1 to a.NAVHeader'length loop
         y(k) := a.NAVHeader(i);
         k := k + 1;
      end loop;

      return y;
   end to_DPB_DCube_Header_array32_v2_6;   
   
   function to_DPB_DCube_Header_array32(a: DPB_DCube_Header) return DPB_DCube_Header_array32 is
      variable y: DPB_DCube_Header_array32;
      variable y1: ROIC_DCube_Header_array32;
      variable y2: ROIC_DCube_Footer_array32;
   begin 
      -- No Header section, THE ARRAY CONTAINS ONLY THE PAYLOAD
      -- DPB Section
      y(1) := PROC_HEADER_FRAME & std_logic_vector(to_unsigned(DPB_DCube_Header_array32'length-1, 24)); -- Command Header + payload size
      y(2)(31 downto DUILEN) := (others => '0');
      y(2)(DUILEN-1 downto 0) := std_logic_vector(a.DUI);
      y(3)(31 downto 16) := (others => '0');
      y(3)(15 downto 0) := a.VP30Status.ExtTemp & a.VP30Status.IntTemp;
      y(4) := a.VP30Status.Stat;
      -- ROIC Header Section (skip header word)
      y1 := to_ROIC_DCube_Header_array32(a.ROICHeader);
      for i in 2 to y1'length loop
         y(i+3) := y1(i);
      end loop;
      -- ROIC Footer Section (skip header word)
      y2 := to_ROIC_DCube_Footer_array32(a.ROICFooter);
      for i in 2 to y2'length loop
         y(i+2+y1'length) := y2(i);
      end loop;
      return y;
   end to_DPB_DCube_Header_array32; 
   
   -- pragma translate_off
   function to_DPConfig_array32 (a: DPConfig) return DPConfig_array32 is
      variable y : DPConfig_array32;
      variable  data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 17; -- In 32-bit elements
   begin
      y(1) := x"61" & std_logic_vector(to_unsigned(PayloadSize,24));
      for i in 1 to PayloadSize loop
         case i is
            when 1  => data32_slv := std_logic_vector(resize(a.ZSIZE	   , 32));
            when 2  => data32_slv := std_logic_vector(resize(a.XSIZE	   , 32));
            when 3  => data32_slv := std_logic_vector(resize(a.YSIZE		, 32));
            when 4  => data32_slv := std_logic_vector(resize(a.IMGSIZE  , 32));
            when 5  => data32_slv := std_logic_vector(resize(a.TAGSIZE	, 32));
            when 6  => data32_slv := std_logic_vector(resize(a.SB_Min   , 32));
            when 7  => data32_slv := std_logic_vector(resize(a.SB_Max   , 32));
            when 8  => data32_slv := std_logic_vector(resize(a.SB_Mode  , 32));
            when 9  => data32_slv := std_logic_vector(resize(unsigned(a.Interleave) , 32));
            when 10 => data32_slv := std_logic_vector(resize(unsigned(a.Mode)       , 32));
            when 11 => data32_slv := std_logic_vector(resize(a.AVGSIZE	  , 32));
            when 12 => data32_slv := std_logic_vector(resize(a.DIAGSIZE   , 32));
            when 13 => data32_slv := std_logic_vector(resize(a.BB_Temp    , 32));
            when 14 => data32_slv := std_logic_vector(resize(unsigned(a.Delta_OPD)  , 32));
            when 15 => data32_slv := std_logic_vector(resize(a.Max_Temp   , 32));
            when 16 => data32_slv := std_logic_vector(resize(a.SB_Min_Cal , 32));
            when 17 => data32_slv := std_logic_vector(resize(a.SB_Max_Cal , 32));
            --when 18 => data32_slv := std_logic_vector(resize(a.Lh_Exp     , 32));
            --when 19 => data32_slv := std_logic_vector(resize(a.DLbb_Exp   , 32));
         end case;
         y(i+1) := data32_slv;
      end loop;
      
      return y;
   end to_DPConfig_array32;
   
   function to_DPConfig_array32 (a: DPConfig; MissingImages : integer) return DPConfig_array32 is
      variable y : DPConfig_array32;
      variable  data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSize : integer := 17; -- In 32-bit elements
   begin
      y(1) := x"61" & std_logic_vector(to_unsigned(PayloadSize,24));
      for i in 1 to PayloadSize loop
         case i is
            when 1  => data32_slv := std_logic_vector(resize(a.ZSIZE	   , 32));
            when 2  => data32_slv := std_logic_vector(resize(a.XSIZE	   , 32));
            when 3  => data32_slv := std_logic_vector(resize(a.YSIZE		, 32));
            when 4  => data32_slv := std_logic_vector(resize(a.IMGSIZE  , 32));
            when 5  => data32_slv := std_logic_vector(resize(a.TAGSIZE	, 32));
            when 6  => data32_slv := std_logic_vector(resize(a.SB_Min   , 32));
            when 7  => data32_slv := std_logic_vector(resize(a.SB_Max   , 32));
            when 8  => data32_slv := std_logic_vector(resize(a.SB_Mode  , 32));
            when 9  => data32_slv := std_logic_vector(resize(unsigned(a.Interleave) , 32));
            when 10 => data32_slv := std_logic_vector(resize(unsigned(a.Mode) + to_unsigned(MissingImages*65536,32) , 32));
            when 11 => data32_slv := std_logic_vector(resize(a.AVGSIZE	  , 32));
            when 12 => data32_slv := std_logic_vector(resize(a.DIAGSIZE   , 32));
            when 13 => data32_slv := std_logic_vector(resize(a.BB_Temp    , 32));
            when 14 => data32_slv := std_logic_vector(resize(unsigned(a.Delta_OPD)  , 32));
            when 15 => data32_slv := std_logic_vector(resize(a.Max_Temp   , 32));
            when 16 => data32_slv := std_logic_vector(resize(a.SB_Min_Cal , 32));
            when 17 => data32_slv := std_logic_vector(resize(a.SB_Max_Cal , 32));
            --when 18 => data32_slv := std_logic_vector(resize(a.Lh_Exp     , 32));
            --when 19 => data32_slv := std_logic_vector(resize(a.DLbb_Exp   , 32));
         end case;
         y(i+1) := data32_slv;
      end loop;
      
      return y;
   end to_DPConfig_array32;   
   -- pragma translate_on
   
   -- private RS232 command 62 for configuring pattern generator via RS232
   function to_PatGenConfig (a: patgen_array8; ValidConfig: boolean) return PatGenConfig is
      variable y : PatGenConfig;
      variable data32 : unsigned(31 downto 0);
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSizeInBytes : integer := PatGen_array8'LENGTH-2; -- In 32-bit elements
      constant PayloadSize : integer := PayloadSizeInBytes/4;
   begin
      -- translate_off
      assert a(1) = x"62" report "Wrong header received, expected 0x62" severity ERROR;
      if ValidConfig then
         assert (to_integer(unsigned(a(2))) = PayloadSizeInBytes) report "Wrong payload size received for command 0x62" severity ERROR;
      end if;
      -- translate_on
      
      for i in 1 to PayloadSize loop
         data32_slv := a(i*4-3 + 2) & a(i*4-2 + 2) & a(i*4-1 + 2) & a(i*4 + 2);
         data32 := unsigned(data32_slv);
         
         case i is
            when 1  =>
               y.Trig :=data32_slv(31);
               y.FrameType   := std_logic_vector(resize(data32, 8));
            when 2  => y.XSize       := resize(data32, XLEN);
            when 3  => y.YSize       := resize(data32, YLEN);
            when 4  => y.ZSize       := resize(data32, ZLEN);
            when 5  => y.DiagSize    := resize(data32, DIAGLEN);
            when 6  => y.PayloadSize := resize(data32, PLLEN);
            when 7  => y.TagSize     := resize(data32, TAGLEN);
            when 8  => y.DiagMode    := std_logic_vector(resize(data32, DIAGMODELEN));
         end case;
      end loop;   
      y.ImagePause := to_unsigned(2, y.ImagePause'LENGTH); -- PDU : Not part of RS232 command (yet).
      return y;
   end to_PatGenConfig;
   
   -- translate_off
   function to_patgen_array8 (a: PatGenConfig) return patgen_array8 is
      variable y : patgen_array8;
      variable data32 : unsigned(31 downto 0);
      variable data32_slv : std_logic_vector(31 downto 0);
      constant PayloadSizeInBytes : integer := PatGen_array8'LENGTH-2; -- In 32-bit elements
      constant PayloadSize : integer := PayloadSizeInBytes/4;
   begin
      y(1) := x"62";
      y(2) := std_logic_vector(to_unsigned(PayloadSizeInBytes,8)); -- Payload size
      
      for i in 1 to PayloadSize loop
         case i is
            when 1 =>
               data32(31) := a.trig;
               data32(30 downto 0) := resize(unsigned(a.FrameType), 31);
            when 2 => data32 := resize(a.XSize, 32);
            when 3 => data32 := resize(a.YSize, 32);
            when 4 => data32 := resize(a.ZSize, 32);
            when 5 => data32 := resize(a.DiagSize, 32);
            when 6 => data32 := resize(a.PayloadSize, 32);
            when 7 => data32 := resize(a.TagSize, 32);
            when 8 => data32 := resize(unsigned(a.DiagMode), 32);
         end case;
         data32_slv := std_logic_vector(data32);
         y(i*4-3 + 2) := data32_slv(31 downto 24); -- MSB
         y(i*4-2 + 2) := data32_slv(23 downto 16);
         y(i*4-1 + 2) := data32_slv(15 downto 8);
         y(i*4 + 2)   := data32_slv(7 downto 0);-- LSB
      end loop;
      
      return y;
   end to_patgen_array8;
   -- translate_on
   
end package body DPB_Define;
