---------------------------------------------------------------------------------------------------
--
-- Title       : div_gen_dval
-- Design      : CAMEL
-- Author      : Patrick Dubois
-- Company     : Telops

---------------------------------------------------------------------------------------------------
--
-- Description : This module adds a "Data Valid" signal to a divider generated by the Core Generator
--
---------------------------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity div_gen_dval is
	generic(
		Latency : integer := 24);
	port(
		CLK 			: in 	STD_LOGIC;
		RST			: in	STD_LOGIC;
		DIV_CE 		: in 	STD_LOGIC;
		DIV_RFD 		: in 	STD_LOGIC;
		DIV_IN_DVAL : in 	std_logic;
		DIV_OUT_DVAL: out STD_LOGIC);
end div_gen_dval;


architecture RTL of div_gen_dval is
signal shift_reg : std_logic_vector(Latency-1 downto 0);
begin
	DIV_OUT_DVAL <= shift_reg(Latency-1);
	
	proc : process(CLK, RST)
	begin
		if rising_edge(CLK) then
			if RST = '1' then
				shift_reg <= (others => '0');
			elsif DIV_CE = '1' then																 
				shift_reg(0) <= DIV_RFD and DIV_IN_DVAL;
				shift_reg(Latency-1 downto 1) <= shift_reg(Latency-2 downto 0);					
			end if;
		end if;
	end process;
	
end RTL;	

--component div_gen_dval
--	generic(
--		Latency : integer := 24);
--	port(
--		CLK 			: in 	STD_LOGIC;
--		RST			: in	STD_LOGIC;
--		DIV_CE 		: in 	STD_LOGIC;
--		DIV_RFD 		: in 	STD_LOGIC;
--		DIV_IN_DVAL : in 	std_logic;
--		DIV_OUT_DVAL: out STD_LOGIC);
--end component;
--
--your_instance : div_gen_dval
--generic map (
--	Latency => 24,
--	ClocksPerDivision => 4)
--port map (
--	CLK => CLK,
--	CLK => RST,
--	DIV_CE => div_Ice,
--	DIV_RFD => div_rfd,
--	DIV_IN_DVAL => div_in_dval,
--	DIV_OUT_DVAL => div_dval);
