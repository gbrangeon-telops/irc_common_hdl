--
--      Project:  Aurora Module Generator version 2.4
--
--         Date:  $Date: 2005/11/07 21:30:52 $
--          Tag:  $Name: i+IP+98818 $
--         File:  $RCSfile: frame_check_vhd.ejava,v $
--          Rev:  $Revision: 1.1.2.4 $
--
--      Company:  Xilinx
-- Contributors:  R. K. Awalt, B. L. Woodard, N. Gulstone, N. Jayarajan
--
--   Disclaimer:  XILINX IS PROVIDING THIS DESIGN, CODE, OR
--                INFORMATION "AS IS" SOLELY FOR USE IN DEVELOPING
--                PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY
--                PROVIDING THIS DESIGN, CODE, OR INFORMATION AS
--                ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE,
--                APPLICATION OR STANDARD, XILINX IS MAKING NO
--                REPRESENTATION THAT THIS IMPLEMENTATION IS FREE
--                FROM ANY CLAIMS OF INFRINGEMENT, AND YOU ARE
--                RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY
--                REQUIRE FOR YOUR IMPLEMENTATION.  XILINX
--                EXPRESSLY DISCLAIMS ANY WARRANTY WHATSOEVER WITH
--                RESPECT TO THE ADEQUACY OF THE IMPLEMENTATION,
--                INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR
--                REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE
--                FROM CLAIMS OF INFRINGEMENT, IMPLIED WARRANTIES
--                OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
--                PURPOSE.
--
--                (c) Copyright 2004 Xilinx, Inc.
--                All rights reserved.
--

--
--  FRAME_CHECK
--
--  Author: Nanditha Jayarajan, Nigel Gulstone
--          Xilinx - Embedded Networking System Engineering Group
--
--
--  Description: This module is a  pattern checker to test the Aurora
--               designs in hardware. The frames generated by FRAME_GEN
--               pass through the Aurora channel and arrive at the frame checker 
--               through the RX User interface. Every time an error is found in
--               the data recieved, the error count is incremented until it 
--               reaches its max value.


library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use WORK.AURORA.all;

-- synthesis translate_off
library UNISIM;
use UNISIM.all;
-- synthesis translate_on


entity FRAME_CHECK is
port
(
    -- User Interface
    RX_D            : in  std_logic_vector(0 to 63); 
    RX_REM          : in  std_logic_vector(0 to 2);     
    RX_SOF_N        : in  std_logic;
    RX_EOF_N        : in  std_logic;
    RX_SRC_RDY_N    : in  std_logic;  

    -- System Interface
    USER_CLK        : in  std_logic;   
    RESET           : in  std_logic;
    ERROR_COUNT     : out std_logic_vector(0 to 7)
  
);
end FRAME_CHECK;



architecture RTL of FRAME_CHECK is

--***********************************Parameter Declarations***************************

    constant DLY : time := 1 ns;

--***************************Internal Register Declarations*************************** 

    signal  in_frame_r          :   std_logic;
    signal  data_r              :   std_logic_vector(0 to 63);
    signal  data_valid_r        :   std_logic;
    signal  error_detected_r    :   std_logic;
    signal  error_count_r       :   std_logic_vector(0 to 8);
    
 
--*********************************Wire Declarations**********************************
   
    signal  data_valid_c        :   std_logic;
    signal  in_frame_c          :   std_logic;
    signal  rem_valid_c         :   std_logic;
    
    signal  error_detected_c    :   std_logic;


begin
--*********************************Main Body of Code**********************************


    --______________________________ Capture incoming data ___________________________    
    --Data is valid when RX_SRC_RDY_N is asserted and data is arriving within a frame
    data_valid_c    <=   in_frame_c and rem_valid_c and not RX_SRC_RDY_N;


    --Data is in a frame if it is a single cycle frame or a multi_cycle frame has started
    in_frame_c      <=   in_frame_r  or  (not RX_SRC_RDY_N and not RX_SOF_N);
    
    
    --Start a multicycle frame when a frame starts without ending on the same cycle. End 
    --the frame when an EOF is detected
    process(USER_CLK)
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(RESET = '1') then   
                in_frame_r  <=  '0' after DLY;
            elsif( (not in_frame_r and not RX_SOF_N and not RX_SRC_RDY_N and RX_EOF_N)='1' ) then
                in_frame_r  <=  '1' after DLY;
            elsif( (in_frame_r and not RX_SRC_RDY_N and not RX_EOF_N)='1' ) then
                in_frame_r  <=  '0' after DLY;
            end if;
        end if;
    end process;
      
      
    --We expect rem to indicate a full word of data on the EOF cycle
    rem_valid_c <=   RX_EOF_N or std_bool(RX_REM = "111");
                


    --Capture valid incoming data, right shifted 1 bit for comparison with the next valid
    --incoming data
    process(USER_CLK)
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(data_valid_c = '1') then
                data_r  <=  (RX_D(63) & RX_D(0 to 62)) after DLY;
            end if;
        end if;
    end process;
 

    --Data in the data register is valid only if it was valid when captured and had no error
    process(USER_CLK)
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(RESET = '1') then
                data_valid_r    <=  '0' after DLY;
            else
                data_valid_r    <=  data_valid_c and not error_detected_c after DLY;
            end if;
        end if;
    end process;


    
    --___________________________ Check incoming data for errors __________________________
         
    
    --An error is detected when valid data from the data register, when right shifted, does not match valid data
    --from the Aurora RX port
    error_detected_c    <=   data_valid_c and data_valid_r and std_bool(RX_D /= data_r);   
    
    
    --We register the error_detected signal for use with the error counter logic
    process(USER_CLK)
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(RESET = '1') then
                error_detected_r    <=  '0' after DLY;
            else
                error_detected_r    <=  error_detected_c after DLY;
            end if;
        end if;
    end process;
    
    
    --We count the total number of errors we detect. By keeping a count we make it less likely that we will miss
    --errors we did not directly observe. This counter must be reset when it reaches its max value
    process(USER_CLK)
    begin
        if(USER_CLK'event and USER_CLK = '1') then
            if(RESET = '1') then
                error_count_r   <=  "000000000" after DLY;
            elsif( (error_detected_r and not error_count_r(0))='1' ) then
                error_count_r   <=  error_count_r + 1 after DLY;
            end if;
        end if;
    end process;            
    
    
    --Here we connect the lower 8 bits of the count (the MSbit is used only to check when the counter reaches
    --max value) to the module output
    ERROR_COUNT <=   error_count_r(1 to 8);    


end RTL;
